module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01662_;
 wire _01664_;
 wire _01665_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01677_;
 wire net3471;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire net3468;
 wire _01693_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01707_;
 wire _01708_;
 wire _01710_;
 wire _01711_;
 wire _01713_;
 wire net3466;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01761_;
 wire _01762_;
 wire _01764_;
 wire _01765_;
 wire clknet_leaf_83_clk_i_regs;
 wire _01767_;
 wire _01768_;
 wire net3477;
 wire _01771_;
 wire net3464;
 wire _01773_;
 wire net3463;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01780_;
 wire _01781_;
 wire _01783_;
 wire _01784_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01815_;
 wire _01816_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire clknet_leaf_84_clk_i_regs;
 wire _01830_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01867_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire net3462;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire net3461;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire net3460;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire net3458;
 wire _02008_;
 wire _02009_;
 wire _02012_;
 wire _02013_;
 wire _02015_;
 wire _02016_;
 wire net3465;
 wire _02019_;
 wire _02020_;
 wire _02022_;
 wire _02023_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02063_;
 wire _02064_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire net3459;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02129_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire clknet_leaf_85_clk_i_regs;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire clknet_leaf_86_clk_i_regs;
 wire _02153_;
 wire _02156_;
 wire _02160_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02171_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02186_;
 wire _02187_;
 wire _02189_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire clknet_leaf_88_clk_i_regs;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02242_;
 wire _02243_;
 wire _02245_;
 wire _02246_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02299_;
 wire _02301_;
 wire _02302_;
 wire _02304_;
 wire _02305_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02322_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02426_;
 wire _02427_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02505_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02853_;
 wire _02855_;
 wire _02856_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire clknet_leaf_92_clk_i_regs;
 wire _02966_;
 wire net3723;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02995_;
 wire net3745;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire net3446;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire net3741;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire net3448;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire net3445;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire net3447;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire clknet_0_clk_i_regs;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire clknet_3_2__leaf_clk_i_regs;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire net3444;
 wire _03280_;
 wire net3744;
 wire clknet_3_7__leaf_clk_i_regs;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire net3449;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire net3432;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire net3442;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03410_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire net3431;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire net3430;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire net3433;
 wire clknet_leaf_2_clk;
 wire _03470_;
 wire _03471_;
 wire clknet_leaf_3_clk;
 wire _03473_;
 wire _03474_;
 wire clknet_leaf_4_clk;
 wire _03476_;
 wire _03477_;
 wire net3427;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire clknet_leaf_6_clk;
 wire _03486_;
 wire net3434;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire net3435;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire net3424;
 wire clknet_leaf_8_clk;
 wire _03546_;
 wire _03547_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire clknet_leaf_9_clk;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire net3422;
 wire net3421;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire net3417;
 wire net3418;
 wire _03697_;
 wire net3429;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire net3415;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire net3419;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire net3412;
 wire _03803_;
 wire net3414;
 wire _03805_;
 wire net3416;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire net3409;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire net3408;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire net3407;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire net3406;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_7_clk;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire net3425;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04038_;
 wire _04039_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04462_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04492_;
 wire _04495_;
 wire _04496_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04656_;
 wire net3440;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire net3746;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire clknet_3_3__leaf_clk_i_regs;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire net3953;
 wire _04734_;
 wire net3952;
 wire net3947;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire net3951;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire net3413;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire net3420;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire net3423;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire net3426;
 wire clknet_leaf_11_clk;
 wire net3405;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire clknet_3_4__leaf_clk_i_regs;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire clknet_leaf_5_clk;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire net3428;
 wire _05082_;
 wire _05083_;
 wire net3404;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire clknet_leaf_1_clk;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire clknet_leaf_0_clk;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire clknet_3_5__leaf_clk_i_regs;
 wire clknet_leaf_12_clk;
 wire _05118_;
 wire clknet_leaf_13_clk;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire net3441;
 wire net3747;
 wire clknet_leaf_26_clk;
 wire _05127_;
 wire _05128_;
 wire net3950;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire net3643;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire net3948;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire net3949;
 wire _05167_;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_27_clk;
 wire _05171_;
 wire _05172_;
 wire clknet_leaf_22_clk;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire clknet_leaf_28_clk;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire clknet_leaf_29_clk;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_21_clk;
 wire _05212_;
 wire _05213_;
 wire clknet_leaf_30_clk;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire clknet_3_0__leaf_clk_i_regs;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire net3871;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire net3402;
 wire net3872;
 wire net3955;
 wire _05253_;
 wire _05254_;
 wire clknet_leaf_13_clk_i_regs;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire clknet_leaf_10_clk_i_regs;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire net3966;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire clknet_leaf_11_clk_i_regs;
 wire net251;
 wire clknet_leaf_12_clk_i_regs;
 wire _05294_;
 wire _05295_;
 wire clknet_leaf_20_clk_i_regs;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire net3931;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire net3969;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire net3963;
 wire clknet_leaf_21_clk_i_regs;
 wire net3921;
 wire _05334_;
 wire _05335_;
 wire net3922;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire clknet_leaf_24_clk;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire clknet_leaf_34_clk;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire net3410;
 wire _05376_;
 wire _05377_;
 wire net3906;
 wire _05379_;
 wire net3907;
 wire clknet_leaf_19_clk;
 wire net3932;
 wire _05383_;
 wire clknet_leaf_15_clk;
 wire _05385_;
 wire net3933;
 wire net3967;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire net3937;
 wire _05395_;
 wire net3964;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire clknet_leaf_16_clk;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire clknet_leaf_35_clk;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire clknet_leaf_36_clk;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_14_clk;
 wire _05433_;
 wire _05434_;
 wire clknet_3_6__leaf_clk_i_regs;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire net3940;
 wire _05441_;
 wire _05442_;
 wire net253;
 wire _05444_;
 wire net3403;
 wire net3912;
 wire _05447_;
 wire net3826;
 wire _05449_;
 wire net3873;
 wire _05451_;
 wire net3934;
 wire _05453_;
 wire net254;
 wire net3900;
 wire _05456_;
 wire net3970;
 wire _05458_;
 wire net3817;
 wire _05460_;
 wire net3773;
 wire _05462_;
 wire _05463_;
 wire net3764;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire net3766;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire net3760;
 wire _05475_;
 wire net3762;
 wire _05477_;
 wire net3751;
 wire net3753;
 wire _05480_;
 wire net3777;
 wire _05482_;
 wire net3736;
 wire _05484_;
 wire net3767;
 wire _05486_;
 wire net3731;
 wire _05488_;
 wire net3792;
 wire _05490_;
 wire net3687;
 wire _05492_;
 wire _05493_;
 wire net3669;
 wire _05495_;
 wire net3674;
 wire _05497_;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_89_clk_i_regs;
 wire net3633;
 wire _05501_;
 wire _05502_;
 wire net3617;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire net3630;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire net3496;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire clknet_leaf_47_clk;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire clknet_leaf_48_clk;
 wire net259;
 wire clknet_leaf_36_clk_i_regs;
 wire _05545_;
 wire _05546_;
 wire net296;
 wire _05548_;
 wire net297;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire clknet_leaf_40_clk_i_regs;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire net433;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire net467;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05586_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire clknet_3_1__leaf_clk_i_regs;
 wire _05594_;
 wire _05595_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05641_;
 wire _05642_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05686_;
 wire _05687_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05728_;
 wire _05729_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05815_;
 wire _05816_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05825_;
 wire _05826_;
 wire _05828_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05867_;
 wire _05868_;
 wire _05870_;
 wire _05872_;
 wire _05874_;
 wire _05876_;
 wire _05878_;
 wire _05880_;
 wire _05881_;
 wire _05884_;
 wire _05886_;
 wire _05888_;
 wire _05890_;
 wire _05893_;
 wire _05895_;
 wire _05897_;
 wire _05899_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05911_;
 wire _05913_;
 wire _05916_;
 wire _05918_;
 wire _05920_;
 wire _05922_;
 wire _05924_;
 wire _05925_;
 wire _05927_;
 wire _05928_;
 wire _05930_;
 wire _05932_;
 wire _05936_;
 wire _05937_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05981_;
 wire _05982_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06025_;
 wire _06026_;
 wire _06028_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06071_;
 wire _06072_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06116_;
 wire _06117_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire net149;
 wire net148;
 wire net147;
 wire _06160_;
 wire _06161_;
 wire net146;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire net145;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire net144;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire net143;
 wire net142;
 wire net141;
 wire _06202_;
 wire _06203_;
 wire net140;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire net139;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire net138;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire net137;
 wire net136;
 wire net135;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire net134;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire net133;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire net132;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire net131;
 wire net130;
 wire net129;
 wire _06288_;
 wire _06289_;
 wire net128;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire net127;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire net126;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire net125;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire net124;
 wire net123;
 wire net122;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire net121;
 wire _06386_;
 wire net120;
 wire _06388_;
 wire _06389_;
 wire net119;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire net118;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire net117;
 wire _06412_;
 wire _06413_;
 wire net116;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire net115;
 wire net114;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire net113;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire net112;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire net111;
 wire _06460_;
 wire _06461_;
 wire net110;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire net109;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire net108;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire net107;
 wire net106;
 wire _06506_;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire net101;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire net100;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire net99;
 wire _06527_;
 wire _06528_;
 wire net98;
 wire net97;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire net96;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire net95;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire net94;
 wire _06553_;
 wire net93;
 wire net92;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire net91;
 wire net90;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire net89;
 wire net88;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire net87;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire net86;
 wire _06595_;
 wire _06596_;
 wire net85;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire net84;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire net83;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire net82;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire net81;
 wire net80;
 wire _07002_;
 wire net79;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire net78;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire net77;
 wire _07044_;
 wire _07045_;
 wire net76;
 wire _07047_;
 wire net75;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire net74;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire net73;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire net72;
 wire _07086_;
 wire _07087_;
 wire net71;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire net70;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire net69;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire net68;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire net67;
 wire _07143_;
 wire net66;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire net65;
 wire _07150_;
 wire _07151_;
 wire net64;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire net63;
 wire net62;
 wire _07163_;
 wire net61;
 wire net60;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire net59;
 wire net58;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire net57;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire net56;
 wire _07181_;
 wire net55;
 wire _07183_;
 wire _07184_;
 wire net54;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire net53;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire net52;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire net51;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire net50;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire net49;
 wire net48;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire net47;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire net46;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire net45;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire net44;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire net43;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire net42;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire net41;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire net40;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire net39;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire net38;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire net37;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire net36;
 wire net35;
 wire net34;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire net33;
 wire _07814_;
 wire _07815_;
 wire net32;
 wire net31;
 wire _07818_;
 wire _07819_;
 wire net30;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire net3918;
 wire net3646;
 wire net3919;
 wire net3832;
 wire _07850_;
 wire net3824;
 wire _07852_;
 wire net3944;
 wire net3865;
 wire net3644;
 wire _07856_;
 wire _07857_;
 wire net3845;
 wire net3855;
 wire clknet_leaf_16_clk_i_regs;
 wire net3748;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire net3856;
 wire _07866_;
 wire net3946;
 wire net3822;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire net3443;
 wire _07874_;
 wire net3638;
 wire net3722;
 wire net3655;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire net3637;
 wire clknet_leaf_91_clk_i_regs;
 wire _07891_;
 wire _07892_;
 wire net3653;
 wire _07894_;
 wire _07895_;
 wire net3652;
 wire _07897_;
 wire net3651;
 wire net3545;
 wire _07900_;
 wire clknet_leaf_90_clk_i_regs;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire net3635;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire net3544;
 wire net3450;
 wire net3632;
 wire net3631;
 wire net3451;
 wire net3627;
 wire net3626;
 wire net3625;
 wire net3624;
 wire net3623;
 wire _07924_;
 wire _07925_;
 wire net3622;
 wire _07927_;
 wire net3621;
 wire net3620;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire net3619;
 wire net3618;
 wire _07935_;
 wire net3634;
 wire net3616;
 wire net3641;
 wire net3614;
 wire _07940_;
 wire _07941_;
 wire net3612;
 wire net3615;
 wire _07944_;
 wire _07945_;
 wire net3453;
 wire net3452;
 wire net3457;
 wire net3454;
 wire _07950_;
 wire _07951_;
 wire net3455;
 wire net3456;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire net3467;
 wire _07960_;
 wire net3469;
 wire _07962_;
 wire net420;
 wire clknet_leaf_80_clk_i_regs;
 wire net3536;
 wire net3481;
 wire net3482;
 wire _07968_;
 wire _07969_;
 wire net3483;
 wire net3484;
 wire net3485;
 wire _07973_;
 wire _07974_;
 wire net3486;
 wire _07976_;
 wire net3488;
 wire net3490;
 wire clknet_leaf_75_clk_i_regs;
 wire _07980_;
 wire net3642;
 wire _07982_;
 wire _07983_;
 wire net3608;
 wire net3513;
 wire _07986_;
 wire _07987_;
 wire net3495;
 wire clknet_leaf_74_clk_i_regs;
 wire clknet_leaf_73_clk_i_regs;
 wire net3497;
 wire _07992_;
 wire _07993_;
 wire net3606;
 wire net3610;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire clknet_leaf_71_clk_i_regs;
 wire net3511;
 wire _08003_;
 wire net3501;
 wire _08005_;
 wire _08006_;
 wire net3503;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire net3507;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire net3508;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire clknet_leaf_67_clk_i_regs;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire net3509;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire clknet_leaf_66_clk_i_regs;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire clknet_leaf_65_clk_i_regs;
 wire clknet_leaf_63_clk_i_regs;
 wire net3516;
 wire net3517;
 wire net3518;
 wire clknet_leaf_61_clk_i_regs;
 wire clknet_leaf_60_clk_i_regs;
 wire net3534;
 wire net3520;
 wire _08105_;
 wire clknet_leaf_57_clk_i_regs;
 wire clknet_leaf_58_clk_i_regs;
 wire net3522;
 wire _08109_;
 wire net3529;
 wire _08111_;
 wire net3530;
 wire _08113_;
 wire clknet_leaf_52_clk_i_regs;
 wire clknet_leaf_51_clk_i_regs;
 wire clknet_leaf_50_clk_i_regs;
 wire net3533;
 wire _08118_;
 wire _08119_;
 wire net3537;
 wire _08121_;
 wire clknet_leaf_48_clk_i_regs;
 wire clknet_leaf_45_clk_i_regs;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire net3543;
 wire clknet_leaf_44_clk_i_regs;
 wire net3546;
 wire net3547;
 wire net3549;
 wire _08132_;
 wire net3550;
 wire _08134_;
 wire _08135_;
 wire net3551;
 wire _08137_;
 wire net3552;
 wire _08139_;
 wire net3557;
 wire net3559;
 wire net3560;
 wire clknet_leaf_39_clk_i_regs;
 wire _08144_;
 wire net3563;
 wire _08146_;
 wire _08147_;
 wire net3565;
 wire net3568;
 wire clknet_leaf_37_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire _08152_;
 wire clknet_leaf_34_clk_i_regs;
 wire net3570;
 wire net3573;
 wire clknet_leaf_29_clk_i_regs;
 wire _08157_;
 wire _08158_;
 wire net3572;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire net3574;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire net3609;
 wire _08171_;
 wire _08172_;
 wire clknet_leaf_27_clk_i_regs;
 wire _08174_;
 wire clknet_leaf_26_clk_i_regs;
 wire net3577;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire net3875;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire net3578;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire net3972;
 wire net3602;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire clknet_leaf_24_clk_i_regs;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire net3888;
 wire net3598;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire net3596;
 wire _08223_;
 wire _08224_;
 wire net3973;
 wire net3594;
 wire _08227_;
 wire _08228_;
 wire net3920;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire net3595;
 wire net3597;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire net3599;
 wire _08244_;
 wire net3929;
 wire net3600;
 wire net3601;
 wire net3874;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire net3579;
 wire net3591;
 wire _08253_;
 wire _08254_;
 wire clknet_leaf_1_clk_i_regs;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire clknet_leaf_2_clk_i_regs;
 wire _08260_;
 wire _08261_;
 wire net3583;
 wire _08263_;
 wire clknet_leaf_17_clk_i_regs;
 wire _08265_;
 wire _08266_;
 wire clknet_leaf_3_clk_i_regs;
 wire _08268_;
 wire clknet_leaf_4_clk_i_regs;
 wire net3585;
 wire clknet_leaf_18_clk_i_regs;
 wire net3957;
 wire net3960;
 wire _08274_;
 wire _08275_;
 wire net3961;
 wire net3956;
 wire _08278_;
 wire _08279_;
 wire net3962;
 wire _08281_;
 wire _08282_;
 wire net3936;
 wire net3930;
 wire net3587;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire net3590;
 wire net3589;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire net3917;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire net3593;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire net3592;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire net3889;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire net3890;
 wire net3891;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire net3603;
 wire net3604;
 wire net3605;
 wire _08352_;
 wire net3607;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire net3613;
 wire _08361_;
 wire net3628;
 wire _08363_;
 wire net3629;
 wire _08365_;
 wire net3881;
 wire _08367_;
 wire net3892;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire net3893;
 wire net3958;
 wire net3894;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire net3636;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire net3895;
 wire _08388_;
 wire _08389_;
 wire net3648;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire clknet_leaf_22_clk_i_regs;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire net3645;
 wire net3639;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire net3640;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire net3866;
 wire net3867;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire net3861;
 wire net3654;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire net3657;
 wire _08457_;
 wire net3800;
 wire net3803;
 wire _08460_;
 wire net3795;
 wire net3807;
 wire net3661;
 wire _08464_;
 wire _08465_;
 wire net3721;
 wire _08467_;
 wire _08468_;
 wire net3662;
 wire net3666;
 wire net3670;
 wire _08472_;
 wire net3679;
 wire _08474_;
 wire _08475_;
 wire net3673;
 wire _08477_;
 wire _08478_;
 wire net3675;
 wire _08480_;
 wire net3676;
 wire _08482_;
 wire net3690;
 wire _08484_;
 wire clknet_leaf_5_clk_i_regs;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire clknet_leaf_6_clk_i_regs;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire clknet_leaf_7_clk_i_regs;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire clknet_leaf_19_clk_i_regs;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire net3586;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire clknet_leaf_8_clk_i_regs;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire net3584;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire net281;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire net3683;
 wire _08549_;
 wire net3684;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire net3685;
 wire net3688;
 wire net3582;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire net3699;
 wire net3695;
 wire net3779;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire net3700;
 wire net3725;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire net3732;
 wire net3780;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire net3705;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire net3581;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire net3588;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire net3713;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire net3728;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire net3730;
 wire _08779_;
 wire net3733;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire net3735;
 wire _08803_;
 wire _08804_;
 wire net3737;
 wire net3756;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire net3774;
 wire net3750;
 wire _08818_;
 wire net3758;
 wire _08820_;
 wire clknet_leaf_0_clk_i_regs;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire net3759;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire net3763;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire net3765;
 wire _08847_;
 wire net3776;
 wire _08849_;
 wire net3787;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire net3853;
 wire net3851;
 wire _08861_;
 wire net3850;
 wire _08863_;
 wire net3862;
 wire _08865_;
 wire net3883;
 wire _08867_;
 wire net3884;
 wire net3977;
 wire _08870_;
 wire net3978;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire net3896;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire net3913;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire net3914;
 wire _08919_;
 wire net3400;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire net3399;
 wire net3401;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire net3857;
 wire _08991_;
 wire net3878;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire net3439;
 wire net3438;
 wire _08998_;
 wire _08999_;
 wire net3868;
 wire _09001_;
 wire net3437;
 wire net3869;
 wire _09004_;
 wire _09005_;
 wire net3870;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire net3436;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire net3411;
 wire clknet_leaf_37_clk;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire clknet_leaf_38_clk;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire net3879;
 wire net3877;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire net3580;
 wire clknet_leaf_39_clk;
 wire _09103_;
 wire _09104_;
 wire net3876;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire clknet_leaf_40_clk;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire clknet_leaf_41_clk;
 wire _09127_;
 wire clknet_leaf_42_clk;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire clknet_leaf_43_clk;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire clknet_leaf_44_clk;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_46_clk;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire clknet_leaf_49_clk;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire net3576;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire clknet_leaf_28_clk_i_regs;
 wire clknet_leaf_50_clk;
 wire _09281_;
 wire clknet_leaf_51_clk;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire clknet_leaf_52_clk;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire clknet_leaf_53_clk;
 wire _09292_;
 wire clknet_leaf_54_clk;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire clknet_leaf_55_clk;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire clknet_leaf_56_clk;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire clknet_leaf_57_clk;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire clknet_leaf_58_clk;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire clknet_leaf_59_clk;
 wire _09540_;
 wire _09541_;
 wire clknet_leaf_60_clk;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire clknet_leaf_61_clk;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire net3575;
 wire _09677_;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire _09680_;
 wire clknet_leaf_66_clk;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire clknet_leaf_72_clk;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire clknet_leaf_75_clk;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire clknet_leaf_78_clk;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire clknet_leaf_79_clk;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire clknet_leaf_80_clk;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire clknet_leaf_83_clk;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire clknet_0_clk;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire clknet_3_0_0_clk;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire clknet_3_1_0_clk;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire clknet_leaf_30_clk_i_regs;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire clknet_3_2_0_clk;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire clknet_3_3_0_clk;
 wire _10417_;
 wire _10418_;
 wire clknet_3_4_0_clk;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire clknet_3_5_0_clk;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire clknet_3_6_0_clk;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire clknet_3_7_0_clk;
 wire _10495_;
 wire clknet_leaf_31_clk_i_regs;
 wire delaynet_0_core_clock;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire net3611;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire delaynet_1_core_clock;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire delaynet_2_core_clock;
 wire delaynet_3_core_clock;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire delaynet_4_core_clock;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire clknet_leaf_32_clk_i_regs;
 wire _10559_;
 wire _10560_;
 wire net3569;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire net256;
 wire net3571;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire clknet_leaf_33_clk_i_regs;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire net257;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire net258;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire clknet_leaf_35_clk_i_regs;
 wire net3567;
 wire _10630_;
 wire net3566;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire net260;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire net261;
 wire _10664_;
 wire net262;
 wire _10666_;
 wire _10667_;
 wire net263;
 wire net264;
 wire net265;
 wire net3562;
 wire _10672_;
 wire net266;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire net267;
 wire net3561;
 wire _10679_;
 wire net268;
 wire _10681_;
 wire net269;
 wire _10683_;
 wire _10684_;
 wire net3558;
 wire _10686_;
 wire net270;
 wire net271;
 wire net272;
 wire _10690_;
 wire net273;
 wire clknet_leaf_41_clk_i_regs;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire net274;
 wire _10740_;
 wire net275;
 wire net276;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net282;
 wire net283;
 wire _10753_;
 wire net284;
 wire net285;
 wire _10756_;
 wire _10757_;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire net292;
 wire _10769_;
 wire net293;
 wire net295;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire clknet_leaf_42_clk_i_regs;
 wire net3564;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire net299;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire net3556;
 wire net3554;
 wire net300;
 wire net301;
 wire net302;
 wire net3555;
 wire _10833_;
 wire net3553;
 wire net3548;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire net304;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire net306;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire net308;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire net311;
 wire _10898_;
 wire net313;
 wire _10900_;
 wire _10901_;
 wire net314;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire net315;
 wire net316;
 wire net317;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire net318;
 wire _10928_;
 wire net319;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire net320;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire net321;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire net322;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire net323;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire net324;
 wire _10990_;
 wire _10991_;
 wire net325;
 wire _10993_;
 wire net326;
 wire net327;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire net328;
 wire _11004_;
 wire net329;
 wire _11006_;
 wire _11007_;
 wire net330;
 wire _11009_;
 wire _11010_;
 wire net331;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire net332;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire net333;
 wire net334;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire net335;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire net336;
 wire clknet_leaf_46_clk_i_regs;
 wire _11045_;
 wire net337;
 wire net338;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire net339;
 wire clknet_leaf_47_clk_i_regs;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire net3540;
 wire _11059_;
 wire net3542;
 wire _11061_;
 wire net3539;
 wire _11063_;
 wire _11064_;
 wire net3538;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire net3535;
 wire net3541;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire net340;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire clknet_leaf_49_clk_i_regs;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire net341;
 wire _11089_;
 wire net342;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire net343;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire net344;
 wire _11115_;
 wire net345;
 wire _11117_;
 wire _11118_;
 wire net346;
 wire _11120_;
 wire net347;
 wire net348;
 wire net349;
 wire clknet_leaf_53_clk_i_regs;
 wire _11125_;
 wire clknet_leaf_54_clk_i_regs;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire net356;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire net357;
 wire _11147_;
 wire net358;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire net359;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire net360;
 wire net361;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire net362;
 wire net363;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire net364;
 wire _11179_;
 wire net365;
 wire _11181_;
 wire net366;
 wire net367;
 wire net368;
 wire clknet_leaf_56_clk_i_regs;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire net3531;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire net369;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire net3532;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire clknet_leaf_55_clk_i_regs;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire net370;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire net3528;
 wire net371;
 wire net3525;
 wire net3524;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire net373;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire net478;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire net375;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire net376;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire net377;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire net379;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire net3526;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire net380;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire net381;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire net3521;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire net382;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire net372;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire net383;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire net384;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire net385;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire net386;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire net387;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire net388;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire clknet_leaf_59_clk_i_regs;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire net389;
 wire net3527;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire net390;
 wire net391;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire net3523;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire net482;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire net393;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire net394;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire net395;
 wire _11728_;
 wire _11729_;
 wire net396;
 wire _11731_;
 wire _11732_;
 wire net397;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire net3519;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire net398;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire net399;
 wire _11795_;
 wire _11796_;
 wire net400;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire net401;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire net402;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire net403;
 wire net404;
 wire _11897_;
 wire net405;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire net406;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire net407;
 wire net408;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire net409;
 wire net410;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire net411;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire clknet_leaf_62_clk_i_regs;
 wire net3515;
 wire _11933_;
 wire _11934_;
 wire net412;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire net3512;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire net413;
 wire _12012_;
 wire _12013_;
 wire net414;
 wire _12015_;
 wire _12016_;
 wire clknet_leaf_64_clk_i_regs;
 wire net415;
 wire net416;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire net3510;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire net417;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire net418;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire net419;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire net421;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire net422;
 wire net423;
 wire net424;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire net425;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire net426;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire net427;
 wire net428;
 wire net429;
 wire _12207_;
 wire _12208_;
 wire net430;
 wire clknet_leaf_68_clk_i_regs;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire net431;
 wire _12225_;
 wire clknet_leaf_69_clk_i_regs;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire net432;
 wire _12241_;
 wire _12242_;
 wire net3506;
 wire net3505;
 wire net3504;
 wire _12246_;
 wire net3502;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire net434;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire net435;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire net436;
 wire _12278_;
 wire _12279_;
 wire net437;
 wire _12281_;
 wire clknet_leaf_70_clk_i_regs;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire net438;
 wire net439;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire net440;
 wire _12327_;
 wire _12328_;
 wire net441;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire net442;
 wire _12339_;
 wire _12340_;
 wire net443;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire net444;
 wire net445;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire net446;
 wire _12366_;
 wire _12367_;
 wire net447;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire net448;
 wire _12378_;
 wire _12379_;
 wire net449;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire net450;
 wire _12396_;
 wire net451;
 wire net452;
 wire net466;
 wire _12400_;
 wire net3499;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire clknet_leaf_72_clk_i_regs;
 wire _12406_;
 wire net3500;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire net3498;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire net3514;
 wire net3492;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire net468;
 wire net471;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire net3491;
 wire _12452_;
 wire net472;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire net473;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire net474;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire net479;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire net3493;
 wire _12490_;
 wire _12491_;
 wire net480;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire net481;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire net483;
 wire net484;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire net485;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire net486;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12561_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12596_;
 wire _12597_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire net3489;
 wire _12627_;
 wire _12628_;
 wire net3494;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12639_;
 wire _12640_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12655_;
 wire net3487;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire net3480;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire net3479;
 wire _12748_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12757_;
 wire _12760_;
 wire _12761_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12831_;
 wire _12832_;
 wire _12834_;
 wire _12836_;
 wire _12837_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire net3478;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12895_;
 wire _12896_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire clknet_leaf_78_clk_i_regs;
 wire net3476;
 wire _12966_;
 wire net3474;
 wire net3473;
 wire _12970_;
 wire _12971_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12990_;
 wire _12991_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13051_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13060_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13080_;
 wire _13081_;
 wire _13083_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13109_;
 wire _13110_;
 wire _13112_;
 wire _13113_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire clknet_leaf_82_clk_i_regs;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire clknet_leaf_76_clk_i_regs;
 wire clknet_leaf_81_clk_i_regs;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire clknet_leaf_79_clk_i_regs;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire clknet_leaf_77_clk_i_regs;
 wire net3472;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire net3470;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire net29;
 wire clk_i_regs;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net150;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit_q[0] ;
 wire \cs_registers_i.mcountinhibit_q[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[9] ;
 wire \cs_registers_i.mhpmcounter[1856] ;
 wire \cs_registers_i.mhpmcounter[1857] ;
 wire \cs_registers_i.mhpmcounter[1858] ;
 wire \cs_registers_i.mhpmcounter[1859] ;
 wire \cs_registers_i.mhpmcounter[1860] ;
 wire \cs_registers_i.mhpmcounter[1861] ;
 wire \cs_registers_i.mhpmcounter[1862] ;
 wire \cs_registers_i.mhpmcounter[1863] ;
 wire \cs_registers_i.mhpmcounter[1864] ;
 wire \cs_registers_i.mhpmcounter[1865] ;
 wire \cs_registers_i.mhpmcounter[1866] ;
 wire \cs_registers_i.mhpmcounter[1867] ;
 wire \cs_registers_i.mhpmcounter[1868] ;
 wire \cs_registers_i.mhpmcounter[1869] ;
 wire \cs_registers_i.mhpmcounter[1870] ;
 wire \cs_registers_i.mhpmcounter[1871] ;
 wire \cs_registers_i.mhpmcounter[1872] ;
 wire \cs_registers_i.mhpmcounter[1873] ;
 wire \cs_registers_i.mhpmcounter[1874] ;
 wire \cs_registers_i.mhpmcounter[1875] ;
 wire \cs_registers_i.mhpmcounter[1876] ;
 wire \cs_registers_i.mhpmcounter[1877] ;
 wire \cs_registers_i.mhpmcounter[1878] ;
 wire \cs_registers_i.mhpmcounter[1879] ;
 wire \cs_registers_i.mhpmcounter[1880] ;
 wire \cs_registers_i.mhpmcounter[1881] ;
 wire \cs_registers_i.mhpmcounter[1882] ;
 wire \cs_registers_i.mhpmcounter[1883] ;
 wire \cs_registers_i.mhpmcounter[1884] ;
 wire \cs_registers_i.mhpmcounter[1885] ;
 wire \cs_registers_i.mhpmcounter[1886] ;
 wire \cs_registers_i.mhpmcounter[1887] ;
 wire \cs_registers_i.mhpmcounter[1888] ;
 wire \cs_registers_i.mhpmcounter[1889] ;
 wire \cs_registers_i.mhpmcounter[1890] ;
 wire \cs_registers_i.mhpmcounter[1891] ;
 wire \cs_registers_i.mhpmcounter[1892] ;
 wire \cs_registers_i.mhpmcounter[1893] ;
 wire \cs_registers_i.mhpmcounter[1894] ;
 wire \cs_registers_i.mhpmcounter[1895] ;
 wire \cs_registers_i.mhpmcounter[1896] ;
 wire \cs_registers_i.mhpmcounter[1897] ;
 wire \cs_registers_i.mhpmcounter[1898] ;
 wire \cs_registers_i.mhpmcounter[1899] ;
 wire \cs_registers_i.mhpmcounter[1900] ;
 wire \cs_registers_i.mhpmcounter[1901] ;
 wire \cs_registers_i.mhpmcounter[1902] ;
 wire \cs_registers_i.mhpmcounter[1903] ;
 wire \cs_registers_i.mhpmcounter[1904] ;
 wire \cs_registers_i.mhpmcounter[1905] ;
 wire \cs_registers_i.mhpmcounter[1906] ;
 wire \cs_registers_i.mhpmcounter[1907] ;
 wire \cs_registers_i.mhpmcounter[1908] ;
 wire \cs_registers_i.mhpmcounter[1909] ;
 wire \cs_registers_i.mhpmcounter[1910] ;
 wire \cs_registers_i.mhpmcounter[1911] ;
 wire \cs_registers_i.mhpmcounter[1912] ;
 wire \cs_registers_i.mhpmcounter[1913] ;
 wire \cs_registers_i.mhpmcounter[1914] ;
 wire \cs_registers_i.mhpmcounter[1915] ;
 wire \cs_registers_i.mhpmcounter[1916] ;
 wire \cs_registers_i.mhpmcounter[1917] ;
 wire \cs_registers_i.mhpmcounter[1918] ;
 wire \cs_registers_i.mhpmcounter[1919] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mstatus_q[2] ;
 wire \cs_registers_i.mstatus_q[3] ;
 wire \cs_registers_i.mstatus_q[4] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_mode_id_o[0] ;
 wire \cs_registers_i.priv_mode_id_o[1] ;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire \ex_block_i.alu_i.imd_val_q_i[0] ;
 wire \ex_block_i.alu_i.imd_val_q_i[10] ;
 wire \ex_block_i.alu_i.imd_val_q_i[11] ;
 wire \ex_block_i.alu_i.imd_val_q_i[12] ;
 wire \ex_block_i.alu_i.imd_val_q_i[13] ;
 wire \ex_block_i.alu_i.imd_val_q_i[14] ;
 wire \ex_block_i.alu_i.imd_val_q_i[15] ;
 wire \ex_block_i.alu_i.imd_val_q_i[16] ;
 wire \ex_block_i.alu_i.imd_val_q_i[17] ;
 wire \ex_block_i.alu_i.imd_val_q_i[18] ;
 wire \ex_block_i.alu_i.imd_val_q_i[19] ;
 wire \ex_block_i.alu_i.imd_val_q_i[1] ;
 wire \ex_block_i.alu_i.imd_val_q_i[20] ;
 wire \ex_block_i.alu_i.imd_val_q_i[21] ;
 wire \ex_block_i.alu_i.imd_val_q_i[22] ;
 wire \ex_block_i.alu_i.imd_val_q_i[23] ;
 wire \ex_block_i.alu_i.imd_val_q_i[24] ;
 wire \ex_block_i.alu_i.imd_val_q_i[25] ;
 wire \ex_block_i.alu_i.imd_val_q_i[26] ;
 wire \ex_block_i.alu_i.imd_val_q_i[27] ;
 wire \ex_block_i.alu_i.imd_val_q_i[28] ;
 wire \ex_block_i.alu_i.imd_val_q_i[29] ;
 wire \ex_block_i.alu_i.imd_val_q_i[2] ;
 wire \ex_block_i.alu_i.imd_val_q_i[30] ;
 wire \ex_block_i.alu_i.imd_val_q_i[31] ;
 wire \ex_block_i.alu_i.imd_val_q_i[32] ;
 wire \ex_block_i.alu_i.imd_val_q_i[33] ;
 wire \ex_block_i.alu_i.imd_val_q_i[34] ;
 wire \ex_block_i.alu_i.imd_val_q_i[35] ;
 wire \ex_block_i.alu_i.imd_val_q_i[36] ;
 wire \ex_block_i.alu_i.imd_val_q_i[37] ;
 wire \ex_block_i.alu_i.imd_val_q_i[38] ;
 wire \ex_block_i.alu_i.imd_val_q_i[39] ;
 wire \ex_block_i.alu_i.imd_val_q_i[3] ;
 wire \ex_block_i.alu_i.imd_val_q_i[40] ;
 wire \ex_block_i.alu_i.imd_val_q_i[41] ;
 wire \ex_block_i.alu_i.imd_val_q_i[42] ;
 wire \ex_block_i.alu_i.imd_val_q_i[43] ;
 wire \ex_block_i.alu_i.imd_val_q_i[44] ;
 wire \ex_block_i.alu_i.imd_val_q_i[45] ;
 wire \ex_block_i.alu_i.imd_val_q_i[46] ;
 wire \ex_block_i.alu_i.imd_val_q_i[47] ;
 wire \ex_block_i.alu_i.imd_val_q_i[48] ;
 wire \ex_block_i.alu_i.imd_val_q_i[49] ;
 wire \ex_block_i.alu_i.imd_val_q_i[4] ;
 wire \ex_block_i.alu_i.imd_val_q_i[50] ;
 wire \ex_block_i.alu_i.imd_val_q_i[51] ;
 wire \ex_block_i.alu_i.imd_val_q_i[52] ;
 wire \ex_block_i.alu_i.imd_val_q_i[53] ;
 wire \ex_block_i.alu_i.imd_val_q_i[54] ;
 wire \ex_block_i.alu_i.imd_val_q_i[55] ;
 wire \ex_block_i.alu_i.imd_val_q_i[56] ;
 wire \ex_block_i.alu_i.imd_val_q_i[57] ;
 wire \ex_block_i.alu_i.imd_val_q_i[58] ;
 wire \ex_block_i.alu_i.imd_val_q_i[59] ;
 wire \ex_block_i.alu_i.imd_val_q_i[5] ;
 wire \ex_block_i.alu_i.imd_val_q_i[60] ;
 wire \ex_block_i.alu_i.imd_val_q_i[61] ;
 wire \ex_block_i.alu_i.imd_val_q_i[62] ;
 wire \ex_block_i.alu_i.imd_val_q_i[63] ;
 wire \ex_block_i.alu_i.imd_val_q_i[6] ;
 wire \ex_block_i.alu_i.imd_val_q_i[7] ;
 wire \ex_block_i.alu_i.imd_val_q_i[8] ;
 wire \ex_block_i.alu_i.imd_val_q_i[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_i ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_i ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.compressed_decoder_i.illegal_instr_o ;
 wire net294;
 wire \if_stage_i.compressed_decoder_i.instr_i[10] ;
 wire net303;
 wire net312;
 wire net305;
 wire net307;
 wire net309;
 wire net298;
 wire \if_stage_i.compressed_decoder_i.instr_i[2] ;
 wire \if_stage_i.compressed_decoder_i.instr_i[3] ;
 wire net310;
 wire \if_stage_i.compressed_decoder_i.instr_i[5] ;
 wire \if_stage_i.compressed_decoder_i.instr_i[6] ;
 wire \if_stage_i.compressed_decoder_i.instr_i[7] ;
 wire clknet_leaf_43_clk_i_regs;
 wire \if_stage_i.compressed_decoder_i.instr_i[9] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[0] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[10] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[11] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[12] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[13] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[14] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[15] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[16] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[17] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[18] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[19] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[1] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[20] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[21] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[22] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[23] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[24] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[25] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[26] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[27] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[28] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[29] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[2] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[30] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[31] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[3] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[4] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[5] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[6] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[7] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[8] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[9] ;
 wire \if_stage_i.compressed_decoder_i.is_compressed_o ;
 wire \if_stage_i.fetch_err ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[0] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[1] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[2] ;
 wire \load_store_unit_i.rdata_q[3] ;
 wire \load_store_unit_i.rdata_q[4] ;
 wire \load_store_unit_i.rdata_q[5] ;
 wire \load_store_unit_i.rdata_q[6] ;
 wire \load_store_unit_i.rdata_q[7] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net3847;
 wire net3649;
 wire net3647;
 wire clknet_leaf_15_clk_i_regs;
 wire net3650;
 wire net3928;
 wire net3899;
 wire net3925;
 wire net3943;
 wire net3924;
 wire net3858;
 wire net3923;
 wire net3805;
 wire net3898;
 wire net3927;
 wire net3910;
 wire net3897;
 wire net3911;
 wire net3971;
 wire net3663;
 wire net3979;
 wire net3976;
 wire net3975;
 wire net3974;
 wire net3656;
 wire net3916;
 wire net3887;
 wire net3864;
 wire net3863;
 wire net378;
 wire net3659;
 wire net3658;
 wire net3860;
 wire net3844;
 wire net3854;
 wire net3842;
 wire net3660;
 wire net3841;
 wire net3840;
 wire net3843;
 wire net3836;
 wire net3711;
 wire net3839;
 wire net3834;
 wire net3835;
 wire net3680;
 wire net3664;
 wire net3825;
 wire net3821;
 wire net3852;
 wire net3838;
 wire net3827;
 wire net3665;
 wire net3859;
 wire net3671;
 wire net3667;
 wire net3809;
 wire net3668;
 wire net3710;
 wire net3691;
 wire net3678;
 wire net3804;
 wire net3802;
 wire net3810;
 wire net3672;
 wire net3833;
 wire net3677;
 wire net3681;
 wire net3682;
 wire net3823;
 wire net3819;
 wire net3799;
 wire net3831;
 wire net3686;
 wire net3798;
 wire net3797;
 wire net3689;
 wire net3692;
 wire net3796;
 wire net3791;
 wire net3789;
 wire net3786;
 wire net3784;
 wire net3693;
 wire net3698;
 wire net3788;
 wire net3696;
 wire net3703;
 wire net3697;
 wire net3829;
 wire net3709;
 wire net3785;
 wire net3701;
 wire net3783;
 wire net3782;
 wire net3702;
 wire net3704;
 wire net3781;
 wire net3706;
 wire net3707;
 wire net3778;
 wire net3708;
 wire net3712;
 wire net3714;
 wire net3715;
 wire net3720;
 wire net3717;
 wire net3769;
 wire net3719;
 wire net3716;
 wire net3816;
 wire net3718;
 wire net3775;
 wire net3724;
 wire net3749;
 wire net3726;
 wire net3727;
 wire net3734;
 wire net3729;
 wire net3752;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3742;
 wire net3743;
 wire net3761;
 wire net3757;
 wire net3820;
 wire net3768;
 wire net3770;
 wire net3755;
 wire net3754;
 wire net3772;
 wire net3771;
 wire net3794;
 wire net3828;
 wire net3790;
 wire net3793;
 wire net3806;
 wire net3801;
 wire net3808;
 wire net3811;
 wire net3815;
 wire net3812;
 wire net3814;
 wire net3813;
 wire net3849;
 wire net3818;
 wire net3848;
 wire net3830;
 wire net3837;
 wire net3915;
 wire net3885;
 wire clknet_leaf_23_clk_i_regs;
 wire net3882;
 wire net3942;
 wire net3938;
 wire net3901;
 wire net3965;
 wire net3926;
 wire net3846;
 wire net3959;
 wire net3935;
 wire net3939;
 wire net3909;
 wire net3905;
 wire net3904;
 wire net3902;
 wire net3908;
 wire net3903;
 wire net3941;
 wire clknet_leaf_14_clk_i_regs;
 wire net255;
 wire net3968;
 wire net252;
 wire net250;
 wire net3954;
 wire net3945;

 sky130_fd_sc_hd__and4bb_4 _13246_ (.A_N(\id_stage_i.controller_i.instr_i[3] ),
    .B_N(\id_stage_i.controller_i.instr_i[2] ),
    .C(\id_stage_i.controller_i.instr_i[1] ),
    .D(net329),
    .X(_07845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1312 ();
 sky130_fd_sc_hd__nor4_4 _13251_ (.A(net348),
    .B(net3839),
    .C(net3840),
    .D(net3836),
    .Y(_07850_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1311 ();
 sky130_fd_sc_hd__and3b_4 _13253_ (.A_N(net3830),
    .B(net325),
    .C(net286),
    .X(_07852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1308 ();
 sky130_fd_sc_hd__nor3b_1 _13257_ (.A(net3842),
    .B(net3837),
    .C_N(net3843),
    .Y(_07856_));
 sky130_fd_sc_hd__and4_4 _13258_ (.A(net385),
    .B(_07850_),
    .C(_07852_),
    .D(_07856_),
    .X(_07857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1304 ();
 sky130_fd_sc_hd__inv_12 _13263_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Y(_07862_));
 sky130_fd_sc_hd__inv_4 _13264_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07863_));
 sky130_fd_sc_hd__nand2_8 _13265_ (.A(_07862_),
    .B(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1303 ();
 sky130_fd_sc_hd__nand2_2 _13267_ (.A(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .B(_07864_),
    .Y(_07866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1301 ();
 sky130_fd_sc_hd__clkinvlp_4 _13270_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_07869_));
 sky130_fd_sc_hd__nor2b_4 _13271_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B_N(\load_store_unit_i.ls_fsm_cs[0] ),
    .Y(_07870_));
 sky130_fd_sc_hd__or3b_4 _13272_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .C_N(\load_store_unit_i.ls_fsm_cs[2] ),
    .X(_07871_));
 sky130_fd_sc_hd__o31ai_4 _13273_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_07869_),
    .A3(_07870_),
    .B1(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1300 ();
 sky130_fd_sc_hd__nand2b_4 _13275_ (.A_N(net3833),
    .B(net391),
    .Y(_07874_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1297 ();
 sky130_fd_sc_hd__nor2_1 _13279_ (.A(net3830),
    .B(net3935),
    .Y(_07878_));
 sky130_fd_sc_hd__and2b_4 _13280_ (.A_N(\id_stage_i.controller_i.instr_i[6] ),
    .B(net325),
    .X(_07879_));
 sky130_fd_sc_hd__nand2_4 _13281_ (.A(net3821),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__o21ai_2 _13282_ (.A1(_07874_),
    .A2(_07878_),
    .B1(_07880_),
    .Y(_07881_));
 sky130_fd_sc_hd__nand4bb_4 _13283_ (.A_N(\id_stage_i.controller_i.instr_i[2] ),
    .B_N(\id_stage_i.controller_i.instr_i[3] ),
    .C(\id_stage_i.controller_i.instr_i[1] ),
    .D(net329),
    .Y(_07882_));
 sky130_fd_sc_hd__nor2_4 _13284_ (.A(net325),
    .B(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__nand2_8 _13285_ (.A(net307),
    .B(net287),
    .Y(_07884_));
 sky130_fd_sc_hd__nor2b_4 _13286_ (.A(\id_stage_i.id_fsm_q ),
    .B_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_07885_));
 sky130_fd_sc_hd__nor2_4 _13287_ (.A(_07884_),
    .B(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__a21oi_4 _13288_ (.A1(_07883_),
    .A2(_07886_),
    .B1(_07872_),
    .Y(_07887_));
 sky130_fd_sc_hd__and3_4 _13289_ (.A(net3832),
    .B(_07881_),
    .C(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1295 ();
 sky130_fd_sc_hd__and2_4 _13292_ (.A(\id_stage_i.controller_i.instr_i[1] ),
    .B(net329),
    .X(_07891_));
 sky130_fd_sc_hd__and4b_4 _13293_ (.A_N(net306),
    .B(net3838),
    .C(_07891_),
    .D(_07879_),
    .X(_07892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1294 ();
 sky130_fd_sc_hd__a211oi_2 _13295_ (.A1(_07883_),
    .A2(_07886_),
    .B1(_07892_),
    .C1(net3754),
    .Y(_07894_));
 sky130_fd_sc_hd__and4b_4 _13296_ (.A_N(net325),
    .B(\id_stage_i.controller_i.instr_i[2] ),
    .C(net329),
    .D(\id_stage_i.controller_i.instr_i[1] ),
    .X(_07895_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1293 ();
 sky130_fd_sc_hd__or3b_4 _13298_ (.A(net307),
    .B(net286),
    .C_N(\id_stage_i.controller_i.instr_i[3] ),
    .X(_07897_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1291 ();
 sky130_fd_sc_hd__or3b_4 _13301_ (.A(net356),
    .B(net3935),
    .C_N(\id_stage_i.controller_i.instr_i[12] ),
    .X(_07900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1290 ();
 sky130_fd_sc_hd__nor3b_2 _13303_ (.A(net305),
    .B(\id_stage_i.id_fsm_q ),
    .C_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_07902_));
 sky130_fd_sc_hd__o22ai_4 _13304_ (.A1(_07897_),
    .A2(_07900_),
    .B1(_07902_),
    .B2(_07884_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_4 _13305_ (.A(_07895_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__nor3_2 _13306_ (.A(net3830),
    .B(net3834),
    .C(_07882_),
    .Y(_07905_));
 sky130_fd_sc_hd__nor2b_4 _13307_ (.A(net3935),
    .B_N(net286),
    .Y(_07906_));
 sky130_fd_sc_hd__o22ai_2 _13308_ (.A1(_07884_),
    .A2(_07885_),
    .B1(_07897_),
    .B2(_07900_),
    .Y(_07907_));
 sky130_fd_sc_hd__a22oi_2 _13309_ (.A1(_07905_),
    .A2(_07906_),
    .B1(_07907_),
    .B2(_07895_),
    .Y(_07908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1289 ();
 sky130_fd_sc_hd__nand4b_1 _13311_ (.A_N(net306),
    .B(net3838),
    .C(_07891_),
    .D(_07879_),
    .Y(_07910_));
 sky130_fd_sc_hd__a22oi_2 _13312_ (.A1(_07894_),
    .A2(_07904_),
    .B1(_07908_),
    .B2(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__nor3_4 _13313_ (.A(net3754),
    .B(_07888_),
    .C(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1278 ();
 sky130_fd_sc_hd__mux4_2 _13325_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net3887),
    .S1(net3864),
    .X(_07924_));
 sky130_fd_sc_hd__nand2_1 _13326_ (.A(net3852),
    .B(_07924_),
    .Y(_07925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1277 ();
 sky130_fd_sc_hd__clkinv_16 _13328_ (.A(net3854),
    .Y(_07927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1275 ();
 sky130_fd_sc_hd__mux4_2 _13331_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S0(net3887),
    .S1(net3866),
    .X(_07930_));
 sky130_fd_sc_hd__nand2_1 _13332_ (.A(_07927_),
    .B(_07930_),
    .Y(_07931_));
 sky130_fd_sc_hd__and3_4 _13333_ (.A(net3848),
    .B(_07925_),
    .C(_07931_),
    .X(_07932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1273 ();
 sky130_fd_sc_hd__clkinv_16 _13336_ (.A(net3884),
    .Y(_07935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1269 ();
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .S(net3852),
    .X(_07940_));
 sky130_fd_sc_hd__nor2b_4 _13342_ (.A(net3873),
    .B_N(net3857),
    .Y(_07941_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1267 ();
 sky130_fd_sc_hd__a22o_1 _13345_ (.A1(net3874),
    .A2(_07940_),
    .B1(net3815),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .X(_07944_));
 sky130_fd_sc_hd__nand2b_4 _13346_ (.A_N(net3854),
    .B(net3893),
    .Y(_07945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1263 ();
 sky130_fd_sc_hd__mux2i_1 _13351_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net3874),
    .Y(_07950_));
 sky130_fd_sc_hd__nand2_8 _13352_ (.A(net3856),
    .B(net3893),
    .Y(_07951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1261 ();
 sky130_fd_sc_hd__mux2i_1 _13355_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S(net3874),
    .Y(_07954_));
 sky130_fd_sc_hd__inv_16 _13356_ (.A(net3849),
    .Y(_07955_));
 sky130_fd_sc_hd__o221ai_1 _13357_ (.A1(net363),
    .A2(_07950_),
    .B1(_07951_),
    .B2(_07954_),
    .C1(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__a21oi_2 _13358_ (.A1(_07935_),
    .A2(_07944_),
    .B1(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__clkinv_16 _13359_ (.A(net3844),
    .Y(_07958_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1260 ();
 sky130_fd_sc_hd__nor2_4 _13361_ (.A(_07958_),
    .B(net3848),
    .Y(_07960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1259 ();
 sky130_fd_sc_hd__nor2b_4 _13363_ (.A(net3857),
    .B_N(net3893),
    .Y(_07962_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1254 ();
 sky130_fd_sc_hd__mux2i_1 _13369_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S(net3861),
    .Y(_07968_));
 sky130_fd_sc_hd__nor2b_4 _13370_ (.A(net3892),
    .B_N(net256),
    .Y(_07969_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1251 ();
 sky130_fd_sc_hd__mux2i_1 _13374_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .S(net3861),
    .Y(_07973_));
 sky130_fd_sc_hd__a22oi_2 _13375_ (.A1(net3810),
    .A2(_07968_),
    .B1(net3809),
    .B2(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1250 ();
 sky130_fd_sc_hd__nor2_4 _13377_ (.A(net3854),
    .B(net3893),
    .Y(_07976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1247 ();
 sky130_fd_sc_hd__mux2i_1 _13381_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .S(net3861),
    .Y(_07980_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1246 ();
 sky130_fd_sc_hd__mux2i_1 _13383_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S(net3861),
    .Y(_07982_));
 sky130_fd_sc_hd__and2_4 _13384_ (.A(net341),
    .B(net256),
    .X(_07983_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1244 ();
 sky130_fd_sc_hd__a22oi_2 _13387_ (.A1(net3804),
    .A2(_07980_),
    .B1(_07982_),
    .B2(net3803),
    .Y(_07986_));
 sky130_fd_sc_hd__and3b_4 _13388_ (.A_N(net3850),
    .B(net3848),
    .C(net3844),
    .X(_07987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1240 ();
 sky130_fd_sc_hd__mux4_2 _13393_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S0(net3882),
    .S1(net3861),
    .X(_07992_));
 sky130_fd_sc_hd__and3_4 _13394_ (.A(net3844),
    .B(net3848),
    .C(net3854),
    .X(_07993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1238 ();
 sky130_fd_sc_hd__mux4_2 _13397_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net3882),
    .S1(net3861),
    .X(_07996_));
 sky130_fd_sc_hd__a22o_4 _13398_ (.A1(net3800),
    .A2(_07992_),
    .B1(net3799),
    .B2(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__a31oi_4 _13399_ (.A1(net3751),
    .A2(_07974_),
    .A3(_07986_),
    .B1(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__o31ai_4 _13400_ (.A1(net3844),
    .A2(_07932_),
    .A3(_07957_),
    .B1(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__a22o_4 _13401_ (.A1(net3842),
    .A2(net3667),
    .B1(net3727),
    .B2(net3728),
    .X(_08000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1236 ();
 sky130_fd_sc_hd__nor2_4 _13404_ (.A(net3941),
    .B(net3935),
    .Y(_08003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1235 ();
 sky130_fd_sc_hd__nor2_4 _13406_ (.A(net3830),
    .B(net286),
    .Y(_08005_));
 sky130_fd_sc_hd__and3_4 _13407_ (.A(net3833),
    .B(net386),
    .C(_08005_),
    .X(_08006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1234 ();
 sky130_fd_sc_hd__clkinv_8 _13409_ (.A(net297),
    .Y(_08008_));
 sky130_fd_sc_hd__clkinv_16 _13410_ (.A(net3935),
    .Y(_08009_));
 sky130_fd_sc_hd__nor2_4 _13411_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__o21ai_0 _13412_ (.A1(net3939),
    .A2(_07850_),
    .B1(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_1 _13413_ (.A(_08006_),
    .B(_08011_),
    .Y(_08012_));
 sky130_fd_sc_hd__inv_2 _13414_ (.A(\id_stage_i.controller_i.instr_i[25] ),
    .Y(_08013_));
 sky130_fd_sc_hd__nor2b_4 _13415_ (.A(net298),
    .B_N(net3935),
    .Y(_08014_));
 sky130_fd_sc_hd__or4_4 _13416_ (.A(\id_stage_i.controller_i.instr_i[27] ),
    .B(\id_stage_i.controller_i.instr_i[29] ),
    .C(\id_stage_i.controller_i.instr_i[28] ),
    .D(\id_stage_i.controller_i.instr_i[31] ),
    .X(_08015_));
 sky130_fd_sc_hd__a21oi_2 _13417_ (.A1(_08013_),
    .A2(_08014_),
    .B1(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nor3b_1 _13418_ (.A(net3935),
    .B(net3843),
    .C_N(net298),
    .Y(_08017_));
 sky130_fd_sc_hd__o21ai_0 _13419_ (.A1(net355),
    .A2(_08017_),
    .B1(net3939),
    .Y(_08018_));
 sky130_fd_sc_hd__nor2b_2 _13420_ (.A(net3935),
    .B_N(net298),
    .Y(_08019_));
 sky130_fd_sc_hd__o21ai_0 _13421_ (.A1(net3843),
    .A2(_08019_),
    .B1(net3837),
    .Y(_08020_));
 sky130_fd_sc_hd__nand3_1 _13422_ (.A(_08016_),
    .B(_08018_),
    .C(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__nor4_2 _13423_ (.A(net3839),
    .B(net367),
    .C(\id_stage_i.controller_i.instr_i[31] ),
    .D(net355),
    .Y(_08022_));
 sky130_fd_sc_hd__nor2_2 _13424_ (.A(\id_stage_i.controller_i.instr_i[25] ),
    .B(net348),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_1 _13425_ (.A(_08022_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__nor2_4 _13426_ (.A(net356),
    .B(net3935),
    .Y(_08025_));
 sky130_fd_sc_hd__a21oi_4 _13427_ (.A1(net3944),
    .A2(_08025_),
    .B1(_08014_),
    .Y(_08026_));
 sky130_fd_sc_hd__nor2_1 _13428_ (.A(_08024_),
    .B(_08026_),
    .Y(_08027_));
 sky130_fd_sc_hd__and2_4 _13429_ (.A(_07845_),
    .B(_07852_),
    .X(_08028_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1233 ();
 sky130_fd_sc_hd__o31ai_4 _13431_ (.A1(net3842),
    .A2(_08021_),
    .A3(_08027_),
    .B1(_08028_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2b_4 _13432_ (.A_N(\id_stage_i.id_fsm_q ),
    .B(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_08031_));
 sky130_fd_sc_hd__nor3_4 _13433_ (.A(_07874_),
    .B(_07884_),
    .C(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__nor2_4 _13434_ (.A(net356),
    .B(_08008_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_1 _13435_ (.A1(net3939),
    .A2(_08014_),
    .B1(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand4b_1 _13436_ (.A_N(net325),
    .B(\id_stage_i.controller_i.instr_i[2] ),
    .C(net329),
    .D(\id_stage_i.controller_i.instr_i[1] ),
    .Y(_08035_));
 sky130_fd_sc_hd__nor3_1 _13437_ (.A(_08035_),
    .B(_07897_),
    .C(_08025_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21oi_1 _13438_ (.A1(_08032_),
    .A2(_08034_),
    .B1(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__inv_4 _13439_ (.A(net286),
    .Y(_08038_));
 sky130_fd_sc_hd__or3_1 _13440_ (.A(net306),
    .B(net339),
    .C(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__and2_4 _13441_ (.A(net307),
    .B(net286),
    .X(_08040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1232 ();
 sky130_fd_sc_hd__nor3b_2 _13443_ (.A(net307),
    .B(net286),
    .C_N(net306),
    .Y(_08042_));
 sky130_fd_sc_hd__o21ai_0 _13444_ (.A1(_08040_),
    .A2(_08042_),
    .B1(net339),
    .Y(_08043_));
 sky130_fd_sc_hd__a21o_4 _13445_ (.A1(_08039_),
    .A2(_08043_),
    .B1(net3834),
    .X(_08044_));
 sky130_fd_sc_hd__nor2b_4 _13446_ (.A(net326),
    .B_N(\id_stage_i.controller_i.instr_i[2] ),
    .Y(_08045_));
 sky130_fd_sc_hd__nor2_2 _13447_ (.A(net306),
    .B(net3830),
    .Y(_08046_));
 sky130_fd_sc_hd__nand2b_4 _13448_ (.A_N(_08045_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand2_8 _13449_ (.A(net334),
    .B(net329),
    .Y(_08048_));
 sky130_fd_sc_hd__a21oi_2 _13450_ (.A1(_08044_),
    .A2(_08047_),
    .B1(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__o2111a_4 _13451_ (.A1(_08003_),
    .A2(_08012_),
    .B1(_08049_),
    .C1(_08030_),
    .D1(_08037_),
    .X(_08050_));
 sky130_fd_sc_hd__or4_4 _13452_ (.A(net3833),
    .B(_07882_),
    .C(_07884_),
    .D(_08031_),
    .X(_08051_));
 sky130_fd_sc_hd__nor3_1 _13453_ (.A(net3940),
    .B(_08010_),
    .C(_08003_),
    .Y(_08052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1231 ();
 sky130_fd_sc_hd__clkinvlp_2 _13455_ (.A(\id_stage_i.controller_i.instr_i[30] ),
    .Y(_08054_));
 sky130_fd_sc_hd__nor2_1 _13456_ (.A(net3839),
    .B(net367),
    .Y(_08055_));
 sky130_fd_sc_hd__nor2_2 _13457_ (.A(\id_stage_i.controller_i.instr_i[26] ),
    .B(\id_stage_i.controller_i.instr_i[31] ),
    .Y(_08056_));
 sky130_fd_sc_hd__nand4_1 _13458_ (.A(_08055_),
    .B(_08054_),
    .C(_08023_),
    .D(_08056_),
    .Y(_08057_));
 sky130_fd_sc_hd__a21oi_4 _13459_ (.A1(net3832),
    .A2(_08057_),
    .B1(_07880_),
    .Y(_08058_));
 sky130_fd_sc_hd__nand4_1 _13460_ (.A(_08058_),
    .B(net3943),
    .C(net3936),
    .D(net3940),
    .Y(_08059_));
 sky130_fd_sc_hd__or3b_1 _13461_ (.A(net3942),
    .B(net3935),
    .C_N(\id_stage_i.controller_i.instr_i[30] ),
    .X(_08060_));
 sky130_fd_sc_hd__nand3b_1 _13462_ (.A_N(\id_stage_i.controller_i.instr_i[30] ),
    .B(net3935),
    .C(net3942),
    .Y(_08061_));
 sky130_fd_sc_hd__a21oi_1 _13463_ (.A1(_08060_),
    .A2(_08061_),
    .B1(net3939),
    .Y(_08062_));
 sky130_fd_sc_hd__a31oi_4 _13464_ (.A1(net3939),
    .A2(_08008_),
    .A3(_08054_),
    .B1(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__nand4_1 _13465_ (.A(_08028_),
    .B(_08055_),
    .C(_08023_),
    .D(_08056_),
    .Y(_08064_));
 sky130_fd_sc_hd__nand4_1 _13466_ (.A(net3833),
    .B(net3939),
    .C(net391),
    .D(_08005_),
    .Y(_08065_));
 sky130_fd_sc_hd__o41a_1 _13467_ (.A1(net3939),
    .A2(_07874_),
    .A3(_07884_),
    .A4(_08031_),
    .B1(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__nor4b_1 _13468_ (.A(net3830),
    .B(net3832),
    .C(net348),
    .D_N(net298),
    .Y(_08067_));
 sky130_fd_sc_hd__nand4_1 _13469_ (.A(net3834),
    .B(net3821),
    .C(_08022_),
    .D(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1230 ();
 sky130_fd_sc_hd__a211o_4 _13471_ (.A1(_08051_),
    .A2(_08068_),
    .B1(net3939),
    .C1(_08009_),
    .X(_08070_));
 sky130_fd_sc_hd__o221ai_4 _13472_ (.A1(_08063_),
    .A2(_08064_),
    .B1(_08066_),
    .B2(net3942),
    .C1(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand2_1 _13473_ (.A(_07845_),
    .B(_07852_),
    .Y(_08072_));
 sky130_fd_sc_hd__o2111ai_1 _13474_ (.A1(net3935),
    .A2(_08054_),
    .B1(_08055_),
    .C1(_08023_),
    .D1(_08056_),
    .Y(_08073_));
 sky130_fd_sc_hd__a2bb2o_2 _13475_ (.A1_N(_08072_),
    .A2_N(_08073_),
    .B1(_08006_),
    .B2(_07850_),
    .X(_08074_));
 sky130_fd_sc_hd__or3_4 _13476_ (.A(net356),
    .B(net298),
    .C(net3935),
    .X(_08075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1229 ();
 sky130_fd_sc_hd__nand4_1 _13478_ (.A(net3833),
    .B(net386),
    .C(_08005_),
    .D(_08075_),
    .Y(_08077_));
 sky130_fd_sc_hd__a21oi_1 _13479_ (.A1(_08051_),
    .A2(_08077_),
    .B1(net3935),
    .Y(_08078_));
 sky130_fd_sc_hd__o21ai_2 _13480_ (.A1(_08074_),
    .A2(_08078_),
    .B1(_08033_),
    .Y(_08079_));
 sky130_fd_sc_hd__o2111a_4 _13481_ (.A1(_08051_),
    .A2(_08052_),
    .B1(_08059_),
    .C1(_08071_),
    .D1(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__or2_4 _13482_ (.A(net3830),
    .B(net286),
    .X(_08081_));
 sky130_fd_sc_hd__nor3b_1 _13483_ (.A(net3835),
    .B(net3838),
    .C_N(net326),
    .Y(_08082_));
 sky130_fd_sc_hd__a21oi_1 _13484_ (.A1(net3835),
    .A2(_08045_),
    .B1(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__nor4_2 _13485_ (.A(_08048_),
    .B(_08081_),
    .C(_08025_),
    .D(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__nor2_1 _13486_ (.A(_08035_),
    .B(_07897_),
    .Y(_08085_));
 sky130_fd_sc_hd__a211o_1 _13487_ (.A1(_08015_),
    .A2(_08033_),
    .B1(_08009_),
    .C1(_08085_),
    .X(_08086_));
 sky130_fd_sc_hd__a221oi_4 _13488_ (.A1(_08044_),
    .A2(_08047_),
    .B1(_08084_),
    .B2(_08086_),
    .C1(_08048_),
    .Y(_08087_));
 sky130_fd_sc_hd__nand2_4 _13489_ (.A(net3939),
    .B(_08009_),
    .Y(_08088_));
 sky130_fd_sc_hd__nor3_1 _13490_ (.A(net3944),
    .B(_08024_),
    .C(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__and2_0 _13491_ (.A(_08022_),
    .B(_08023_),
    .X(_08090_));
 sky130_fd_sc_hd__a32oi_1 _13492_ (.A1(_08016_),
    .A2(_08018_),
    .A3(_08020_),
    .B1(_08014_),
    .B2(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__o31ai_2 _13493_ (.A1(net3842),
    .A2(_08091_),
    .A3(_08089_),
    .B1(_08028_),
    .Y(_08092_));
 sky130_fd_sc_hd__nand3_4 _13494_ (.A(_07883_),
    .B(_08040_),
    .C(net3818),
    .Y(_08093_));
 sky130_fd_sc_hd__nand3_4 _13495_ (.A(_08092_),
    .B(_08093_),
    .C(_08087_),
    .Y(_08094_));
 sky130_fd_sc_hd__a21oi_4 _13496_ (.A1(_08080_),
    .A2(_08050_),
    .B1(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1220 ();
 sky130_fd_sc_hd__mux4_2 _13506_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net3923),
    .S1(net3909),
    .X(_08105_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1217 ();
 sky130_fd_sc_hd__clkinv_16 _13510_ (.A(net3902),
    .Y(_08109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1216 ();
 sky130_fd_sc_hd__nor2_4 _13512_ (.A(net3896),
    .B(_08109_),
    .Y(_08111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1215 ();
 sky130_fd_sc_hd__or3_4 _13514_ (.A(net3896),
    .B(net3900),
    .C(net3916),
    .X(_08113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1211 ();
 sky130_fd_sc_hd__mux2i_1 _13519_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .S(net267),
    .Y(_08118_));
 sky130_fd_sc_hd__or3b_4 _13520_ (.A(net3896),
    .B(net3900),
    .C_N(net3913),
    .X(_08119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1210 ();
 sky130_fd_sc_hd__mux2i_1 _13522_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S(net267),
    .Y(_08121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1208 ();
 sky130_fd_sc_hd__o221ai_1 _13525_ (.A1(_08113_),
    .A2(_08118_),
    .B1(_08119_),
    .B2(_08121_),
    .C1(net3898),
    .Y(_08124_));
 sky130_fd_sc_hd__a21oi_1 _13526_ (.A1(_08105_),
    .A2(_08111_),
    .B1(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__and2_4 _13527_ (.A(net3896),
    .B(net3902),
    .X(_08126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1203 ();
 sky130_fd_sc_hd__mux4_2 _13533_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net3920),
    .S1(net3907),
    .X(_08132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1202 ();
 sky130_fd_sc_hd__mux4_2 _13535_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S0(net3920),
    .S1(net3907),
    .X(_08134_));
 sky130_fd_sc_hd__nor2b_4 _13536_ (.A(net3902),
    .B_N(net3896),
    .Y(_08135_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1201 ();
 sky130_fd_sc_hd__a22oi_2 _13538_ (.A1(_08126_),
    .A2(_08132_),
    .B1(_08134_),
    .B2(net3796),
    .Y(_08137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1200 ();
 sky130_fd_sc_hd__nor2b_4 _13540_ (.A(net3913),
    .B_N(net283),
    .Y(_08139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1196 ();
 sky130_fd_sc_hd__mux2i_1 _13545_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .S(net309),
    .Y(_08144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1195 ();
 sky130_fd_sc_hd__mux2i_1 _13547_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S(net309),
    .Y(_08146_));
 sky130_fd_sc_hd__and2_4 _13548_ (.A(net3908),
    .B(net283),
    .X(_08147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1191 ();
 sky130_fd_sc_hd__a221oi_1 _13553_ (.A1(net3793),
    .A2(_08144_),
    .B1(_08146_),
    .B2(net3791),
    .C1(net3896),
    .Y(_08152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1187 ();
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net309),
    .X(_08157_));
 sky130_fd_sc_hd__nor2b_4 _13559_ (.A(net3908),
    .B_N(net3925),
    .Y(_08158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1186 ();
 sky130_fd_sc_hd__or2_4 _13561_ (.A(net3898),
    .B(net3902),
    .X(_08160_));
 sky130_fd_sc_hd__a221o_1 _13562_ (.A1(net3909),
    .A2(_08157_),
    .B1(net3789),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .C1(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__o21ai_0 _13563_ (.A1(net3898),
    .A2(_08152_),
    .B1(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__mux4_2 _13564_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S0(net3920),
    .S1(net3907),
    .X(_08163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1185 ();
 sky130_fd_sc_hd__mux4_2 _13566_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S0(net3920),
    .S1(net3907),
    .X(_08165_));
 sky130_fd_sc_hd__a22oi_2 _13567_ (.A1(_08126_),
    .A2(_08163_),
    .B1(_08165_),
    .B2(net3796),
    .Y(_08166_));
 sky130_fd_sc_hd__a22o_4 _13568_ (.A1(_08125_),
    .A2(_08137_),
    .B1(_08162_),
    .B2(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__inv_6 _13569_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Y(_08168_));
 sky130_fd_sc_hd__clkinv_16 _13570_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Y(_08169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1184 ();
 sky130_fd_sc_hd__nor2_4 _13572_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_08171_));
 sky130_fd_sc_hd__nand3_4 _13573_ (.A(_08168_),
    .B(_08169_),
    .C(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1183 ();
 sky130_fd_sc_hd__nor2_1 _13575_ (.A(net3727),
    .B(_08172_),
    .Y(_08174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1181 ();
 sky130_fd_sc_hd__o22ai_1 _13578_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .B2(net3787),
    .Y(_08177_));
 sky130_fd_sc_hd__a211oi_1 _13579_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_08167_),
    .B1(_08174_),
    .C1(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__o21ai_1 _13580_ (.A1(_08000_),
    .A2(net299),
    .B1(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__xor2_1 _13581_ (.A(_08179_),
    .B(_07866_),
    .X(_08180_));
 sky130_fd_sc_hd__nor3_2 _13582_ (.A(net356),
    .B(net298),
    .C(net3935),
    .Y(_08181_));
 sky130_fd_sc_hd__o21ai_0 _13583_ (.A1(_08081_),
    .A2(_08181_),
    .B1(_07884_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21oi_1 _13584_ (.A1(net330),
    .A2(_08182_),
    .B1(_07886_),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2b_1 _13585_ (.A(net3831),
    .B_N(net3830),
    .Y(_08184_));
 sky130_fd_sc_hd__a2bb2oi_1 _13586_ (.A1_N(net3838),
    .A2_N(_08184_),
    .B1(_08005_),
    .B2(net325),
    .Y(_08185_));
 sky130_fd_sc_hd__o21ai_2 _13587_ (.A1(_08040_),
    .A2(_08042_),
    .B1(_08045_),
    .Y(_08186_));
 sky130_fd_sc_hd__o21ai_2 _13588_ (.A1(net306),
    .A2(_08185_),
    .B1(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__and3_4 _13589_ (.A(net3834),
    .B(_07845_),
    .C(_08040_),
    .X(_08188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1180 ();
 sky130_fd_sc_hd__a222oi_1 _13591_ (.A1(_08038_),
    .A2(_07892_),
    .B1(net3935),
    .B2(_08188_),
    .C1(_07883_),
    .C2(_07886_),
    .Y(_08190_));
 sky130_fd_sc_hd__o2111a_4 _13592_ (.A1(_08035_),
    .A2(_08183_),
    .B1(_08187_),
    .C1(_08190_),
    .D1(_07891_),
    .X(_08191_));
 sky130_fd_sc_hd__nor2_4 _13593_ (.A(_08191_),
    .B(net3754),
    .Y(_08192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1179 ();
 sky130_fd_sc_hd__o31a_1 _13595_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_07869_),
    .A3(_07870_),
    .B1(_07871_),
    .X(_08194_));
 sky130_fd_sc_hd__and3_1 _13596_ (.A(net3938),
    .B(_07895_),
    .C(_08042_),
    .X(_08195_));
 sky130_fd_sc_hd__o22ai_1 _13597_ (.A1(_08188_),
    .A2(_08085_),
    .B1(_08195_),
    .B2(net3935),
    .Y(_08196_));
 sky130_fd_sc_hd__nand4_1 _13598_ (.A(_08194_),
    .B(_07891_),
    .C(_08187_),
    .D(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1177 ();
 sky130_fd_sc_hd__nor2_1 _13601_ (.A(net3723),
    .B(_08167_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21oi_1 _13602_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net3723),
    .B1(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nor3_4 _13603_ (.A(net3754),
    .B(net431),
    .C(net3720),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_1 _13604_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(net3665),
    .Y(_08203_));
 sky130_fd_sc_hd__o21ai_4 _13605_ (.A1(net269),
    .A2(_08201_),
    .B1(_08203_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21o_4 _13606_ (.A1(_08050_),
    .A2(_08080_),
    .B1(_08094_),
    .X(_08205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1176 ();
 sky130_fd_sc_hd__xnor2_1 _13608_ (.A(_08000_),
    .B(_08205_),
    .Y(_08207_));
 sky130_fd_sc_hd__xnor2_1 _13609_ (.A(_08204_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__nor2_1 _13610_ (.A(_08208_),
    .B(net3756),
    .Y(_08209_));
 sky130_fd_sc_hd__a21oi_4 _13611_ (.A1(net3756),
    .A2(_08180_),
    .B1(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1174 ();
 sky130_fd_sc_hd__mux4_2 _13614_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net3884),
    .S1(net3872),
    .X(_08213_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(net295),
    .B(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__mux4_2 _13616_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S0(net3885),
    .S1(net3870),
    .X(_08215_));
 sky130_fd_sc_hd__nand2_1 _13617_ (.A(net3817),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__and3_4 _13618_ (.A(net3848),
    .B(_08214_),
    .C(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .S(net3850),
    .X(_08218_));
 sky130_fd_sc_hd__a22o_4 _13620_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .A2(net3816),
    .B1(_08218_),
    .B2(net3871),
    .X(_08219_));
 sky130_fd_sc_hd__mux2i_1 _13621_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net3871),
    .Y(_08220_));
 sky130_fd_sc_hd__mux2i_1 _13622_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(net3871),
    .Y(_08221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1173 ();
 sky130_fd_sc_hd__o221ai_2 _13624_ (.A1(net3813),
    .A2(_08220_),
    .B1(_08221_),
    .B2(net428),
    .C1(net3812),
    .Y(_08223_));
 sky130_fd_sc_hd__a21oi_4 _13625_ (.A1(_07935_),
    .A2(_08219_),
    .B1(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1171 ();
 sky130_fd_sc_hd__mux2i_1 _13628_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S(net3869),
    .Y(_08227_));
 sky130_fd_sc_hd__mux2i_1 _13629_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .S(net3869),
    .Y(_08228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1170 ();
 sky130_fd_sc_hd__a22oi_1 _13631_ (.A1(net3811),
    .A2(_08227_),
    .B1(_08228_),
    .B2(net3808),
    .Y(_08230_));
 sky130_fd_sc_hd__mux2i_1 _13632_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .S(net3869),
    .Y(_08231_));
 sky130_fd_sc_hd__mux2i_1 _13633_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S(net3869),
    .Y(_08232_));
 sky130_fd_sc_hd__a22oi_2 _13634_ (.A1(net3806),
    .A2(_08231_),
    .B1(_08232_),
    .B2(net3802),
    .Y(_08233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1168 ();
 sky130_fd_sc_hd__mux4_2 _13637_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S0(net3884),
    .S1(net3868),
    .X(_08236_));
 sky130_fd_sc_hd__mux4_2 _13638_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net3884),
    .S1(net3868),
    .X(_08237_));
 sky130_fd_sc_hd__a22o_4 _13639_ (.A1(net3801),
    .A2(_08236_),
    .B1(_08237_),
    .B2(net3798),
    .X(_08238_));
 sky130_fd_sc_hd__a31oi_4 _13640_ (.A1(_08233_),
    .A2(_08230_),
    .A3(net3752),
    .B1(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__o31ai_4 _13641_ (.A1(net3846),
    .A2(_08217_),
    .A3(_08224_),
    .B1(net281),
    .Y(_08240_));
 sky130_fd_sc_hd__a22o_4 _13642_ (.A1(net3843),
    .A2(net3667),
    .B1(_08240_),
    .B2(net3728),
    .X(_08241_));
 sky130_fd_sc_hd__a211oi_4 _13643_ (.A1(_08080_),
    .A2(_08050_),
    .B1(_07857_),
    .C1(_08094_),
    .Y(_08242_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1167 ();
 sky130_fd_sc_hd__nand2_1 _13645_ (.A(_08241_),
    .B(_08242_),
    .Y(_08244_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1159 ();
 sky130_fd_sc_hd__mux4_2 _13654_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net309),
    .S1(net3914),
    .X(_08253_));
 sky130_fd_sc_hd__nand2_1 _13655_ (.A(net3901),
    .B(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1158 ();
 sky130_fd_sc_hd__mux4_2 _13657_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S0(net309),
    .S1(net3914),
    .X(_08256_));
 sky130_fd_sc_hd__nand2_1 _13658_ (.A(_08109_),
    .B(_08256_),
    .Y(_08257_));
 sky130_fd_sc_hd__nor2b_4 _13659_ (.A(net3896),
    .B_N(net3898),
    .Y(_08258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1157 ();
 sky130_fd_sc_hd__nand3_2 _13661_ (.A(_08254_),
    .B(_08257_),
    .C(net3784),
    .Y(_08260_));
 sky130_fd_sc_hd__nand2_8 _13662_ (.A(net3903),
    .B(net3912),
    .Y(_08261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1156 ();
 sky130_fd_sc_hd__mux2_1 _13664_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(net309),
    .X(_08263_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1155 ();
 sky130_fd_sc_hd__mux2_1 _13666_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net309),
    .X(_08265_));
 sky130_fd_sc_hd__nand2b_4 _13667_ (.A_N(net3902),
    .B(net3913),
    .Y(_08266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1154 ();
 sky130_fd_sc_hd__o22ai_2 _13669_ (.A1(net3783),
    .A2(_08263_),
    .B1(_08265_),
    .B2(net3782),
    .Y(_08268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1149 ();
 sky130_fd_sc_hd__mux2_1 _13675_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .S(net439),
    .X(_08274_));
 sky130_fd_sc_hd__and2b_4 _13676_ (.A_N(net3902),
    .B(net3931),
    .X(_08275_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1147 ();
 sky130_fd_sc_hd__a221oi_1 _13679_ (.A1(net3901),
    .A2(_08274_),
    .B1(_08275_),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .C1(net3915),
    .Y(_08278_));
 sky130_fd_sc_hd__nor2_2 _13680_ (.A(net3896),
    .B(net3898),
    .Y(_08279_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1146 ();
 sky130_fd_sc_hd__o21ai_2 _13682_ (.A1(_08268_),
    .A2(_08278_),
    .B1(net3781),
    .Y(_08281_));
 sky130_fd_sc_hd__nor2b_4 _13683_ (.A(net3902),
    .B_N(net3913),
    .Y(_08282_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1143 ();
 sky130_fd_sc_hd__mux2_1 _13687_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S(net3927),
    .X(_08286_));
 sky130_fd_sc_hd__nand2_8 _13688_ (.A(net3896),
    .B(net3899),
    .Y(_08287_));
 sky130_fd_sc_hd__a21oi_1 _13689_ (.A1(net3779),
    .A2(_08286_),
    .B1(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__mux2_1 _13690_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .S(net3927),
    .X(_08289_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S(net3927),
    .X(_08290_));
 sky130_fd_sc_hd__mux2_1 _13692_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .S(net3927),
    .X(_08291_));
 sky130_fd_sc_hd__nor2_4 _13693_ (.A(net3902),
    .B(net3908),
    .Y(_08292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1141 ();
 sky130_fd_sc_hd__a222oi_1 _13696_ (.A1(net266),
    .A2(_08289_),
    .B1(_08290_),
    .B2(net412),
    .C1(_08291_),
    .C2(net3777),
    .Y(_08295_));
 sky130_fd_sc_hd__mux4_2 _13697_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net3927),
    .S1(net3911),
    .X(_08296_));
 sky130_fd_sc_hd__mux4_2 _13698_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S0(net3927),
    .S1(net3911),
    .X(_08297_));
 sky130_fd_sc_hd__mux2i_1 _13699_ (.A0(_08296_),
    .A1(_08297_),
    .S(_08109_),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2b_4 _13700_ (.A(net3898),
    .B_N(net3896),
    .Y(_08299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1140 ();
 sky130_fd_sc_hd__a22oi_2 _13702_ (.A1(_08295_),
    .A2(_08288_),
    .B1(_08298_),
    .B2(net3774),
    .Y(_08301_));
 sky130_fd_sc_hd__nand3_4 _13703_ (.A(_08301_),
    .B(_08281_),
    .C(_08260_),
    .Y(_08302_));
 sky130_fd_sc_hd__o22ai_1 _13704_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .B2(net3787),
    .Y(_08303_));
 sky130_fd_sc_hd__a21oi_1 _13705_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net375),
    .B1(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__o21ai_0 _13706_ (.A1(_08172_),
    .A2(_08240_),
    .B1(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _13707_ (.A(net3756),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__o211ai_1 _13708_ (.A1(net299),
    .A2(_08241_),
    .B1(_08244_),
    .C1(_08306_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand4_1 _13709_ (.A(net385),
    .B(net3820),
    .C(net3819),
    .D(_07852_),
    .Y(_08308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1139 ();
 sky130_fd_sc_hd__nor2_1 _13711_ (.A(net3721),
    .B(net375),
    .Y(_08310_));
 sky130_fd_sc_hd__a21oi_1 _13712_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(net3721),
    .B1(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand2_2 _13713_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(net3665),
    .Y(_08312_));
 sky130_fd_sc_hd__o21ai_4 _13714_ (.A1(net3666),
    .A2(_08311_),
    .B1(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_2 _13715_ (.A(net3744),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__nand2_2 _13716_ (.A(net3820),
    .B(net3819),
    .Y(_08315_));
 sky130_fd_sc_hd__nor3_4 _13717_ (.A(_08038_),
    .B(_07880_),
    .C(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1138 ();
 sky130_fd_sc_hd__nand3_1 _13719_ (.A(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .B(_08316_),
    .C(_07864_),
    .Y(_08318_));
 sky130_fd_sc_hd__nand2_2 _13720_ (.A(_08314_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__xnor2_2 _13721_ (.A(_08307_),
    .B(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__inv_1 _13722_ (.A(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1137 ();
 sky130_fd_sc_hd__mux4_2 _13724_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net3889),
    .S1(net3875),
    .X(_08323_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(net3855),
    .B(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__mux4_2 _13726_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S0(net3889),
    .S1(net3875),
    .X(_08325_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_07927_),
    .B(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__and3_4 _13728_ (.A(net3848),
    .B(_08324_),
    .C(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__mux2_1 _13729_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .S(net3854),
    .X(_08328_));
 sky130_fd_sc_hd__a22o_1 _13730_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .A2(net296),
    .B1(_08328_),
    .B2(net3875),
    .X(_08329_));
 sky130_fd_sc_hd__mux2i_1 _13731_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net3875),
    .Y(_08330_));
 sky130_fd_sc_hd__mux2i_1 _13732_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net3875),
    .Y(_08331_));
 sky130_fd_sc_hd__o221ai_1 _13733_ (.A1(net363),
    .A2(_08330_),
    .B1(_08331_),
    .B2(net426),
    .C1(_07955_),
    .Y(_08332_));
 sky130_fd_sc_hd__a21oi_1 _13734_ (.A1(_07935_),
    .A2(_08329_),
    .B1(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__mux2i_1 _13735_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S(net3875),
    .Y(_08334_));
 sky130_fd_sc_hd__mux2i_1 _13736_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .S(net3875),
    .Y(_08335_));
 sky130_fd_sc_hd__a22oi_1 _13737_ (.A1(net3811),
    .A2(_08334_),
    .B1(_08335_),
    .B2(net3808),
    .Y(_08336_));
 sky130_fd_sc_hd__mux2i_1 _13738_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .S(net3875),
    .Y(_08337_));
 sky130_fd_sc_hd__mux2i_1 _13739_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S(net3875),
    .Y(_08338_));
 sky130_fd_sc_hd__a22oi_1 _13740_ (.A1(net3805),
    .A2(_08337_),
    .B1(_08338_),
    .B2(net3802),
    .Y(_08339_));
 sky130_fd_sc_hd__mux4_2 _13741_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net3890),
    .S1(net3865),
    .X(_08340_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1135 ();
 sky130_fd_sc_hd__mux4_2 _13744_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S0(net3890),
    .S1(net3865),
    .X(_08343_));
 sky130_fd_sc_hd__a22o_4 _13745_ (.A1(net3798),
    .A2(_08340_),
    .B1(_08343_),
    .B2(net275),
    .X(_08344_));
 sky130_fd_sc_hd__a31oi_2 _13746_ (.A1(net3752),
    .A2(_08336_),
    .A3(_08339_),
    .B1(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__o31ai_2 _13747_ (.A1(net3844),
    .A2(_08327_),
    .A3(_08333_),
    .B1(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__nand2_2 _13748_ (.A(_07888_),
    .B(net3719),
    .Y(_08347_));
 sky130_fd_sc_hd__nand3_4 _13749_ (.A(net3832),
    .B(_07881_),
    .C(_07887_),
    .Y(_08348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1132 ();
 sky130_fd_sc_hd__a22o_4 _13753_ (.A1(_07905_),
    .A2(_07906_),
    .B1(_07907_),
    .B2(_07895_),
    .X(_08352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1131 ();
 sky130_fd_sc_hd__o21ai_0 _13755_ (.A1(_07892_),
    .A2(_08352_),
    .B1(net3749),
    .Y(_08354_));
 sky130_fd_sc_hd__a21oi_4 _13756_ (.A1(_07895_),
    .A2(_07903_),
    .B1(net3754),
    .Y(_08355_));
 sky130_fd_sc_hd__a21boi_4 _13757_ (.A1(_07887_),
    .A2(_07908_),
    .B1_N(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__a32o_4 _13758_ (.A1(net285),
    .A2(net3740),
    .A3(_08354_),
    .B1(_08356_),
    .B2(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .X(_08357_));
 sky130_fd_sc_hd__nand2_4 _13759_ (.A(_08348_),
    .B(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__nand2_8 _13760_ (.A(_08347_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1130 ();
 sky130_fd_sc_hd__mux2i_1 _13762_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .S(net3926),
    .Y(_08361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1129 ();
 sky130_fd_sc_hd__mux2i_1 _13764_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net3926),
    .Y(_08363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1128 ();
 sky130_fd_sc_hd__a221oi_1 _13766_ (.A1(net263),
    .A2(_08361_),
    .B1(_08363_),
    .B2(net413),
    .C1(net3896),
    .Y(_08365_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1127 ();
 sky130_fd_sc_hd__mux2_1 _13768_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net346),
    .X(_08367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1126 ();
 sky130_fd_sc_hd__a221o_1 _13770_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .A2(_08158_),
    .B1(_08367_),
    .B2(net3910),
    .C1(_08160_),
    .X(_08369_));
 sky130_fd_sc_hd__o21ai_2 _13771_ (.A1(net3898),
    .A2(_08365_),
    .B1(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__mux4_2 _13772_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net3923),
    .S1(net3910),
    .X(_08371_));
 sky130_fd_sc_hd__mux4_2 _13773_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S0(net3924),
    .S1(net3910),
    .X(_08372_));
 sky130_fd_sc_hd__a22oi_2 _13774_ (.A1(_08126_),
    .A2(_08371_),
    .B1(_08372_),
    .B2(net3796),
    .Y(_08373_));
 sky130_fd_sc_hd__nand2b_4 _13775_ (.A_N(net3908),
    .B(net3903),
    .Y(_08374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1123 ();
 sky130_fd_sc_hd__mux2i_1 _13779_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .S(net3924),
    .Y(_08378_));
 sky130_fd_sc_hd__nor2_1 _13780_ (.A(_08374_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__mux2i_1 _13781_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .S(net3924),
    .Y(_08380_));
 sky130_fd_sc_hd__nor3_1 _13782_ (.A(net3902),
    .B(net3910),
    .C(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__mux2i_1 _13783_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S(net3924),
    .Y(_08382_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1122 ();
 sky130_fd_sc_hd__mux2i_1 _13785_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S(net3924),
    .Y(_08384_));
 sky130_fd_sc_hd__o22ai_1 _13786_ (.A1(_08266_),
    .A2(_08382_),
    .B1(_08384_),
    .B2(_08261_),
    .Y(_08385_));
 sky130_fd_sc_hd__nor4_2 _13787_ (.A(_08287_),
    .B(_08379_),
    .C(_08381_),
    .D(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1121 ();
 sky130_fd_sc_hd__mux4_2 _13789_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S0(net3924),
    .S1(net3910),
    .X(_08388_));
 sky130_fd_sc_hd__or3b_4 _13790_ (.A(net3896),
    .B(net3903),
    .C_N(net3899),
    .X(_08389_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1120 ();
 sky130_fd_sc_hd__nand3b_1 _13792_ (.A_N(net3896),
    .B(net3899),
    .C(net3903),
    .Y(_08391_));
 sky130_fd_sc_hd__mux4_2 _13793_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net3924),
    .S1(net3910),
    .X(_08392_));
 sky130_fd_sc_hd__o22ai_1 _13794_ (.A1(_08388_),
    .A2(_08389_),
    .B1(_08391_),
    .B2(_08392_),
    .Y(_08393_));
 sky130_fd_sc_hd__a211oi_2 _13795_ (.A1(_08370_),
    .A2(_08373_),
    .B1(_08386_),
    .C1(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__nor2_1 _13796_ (.A(_08168_),
    .B(net3716),
    .Y(_08395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1119 ();
 sky130_fd_sc_hd__o22ai_1 _13798_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .B2(net3787),
    .Y(_08397_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_08172_),
    .B(net3719),
    .Y(_08398_));
 sky130_fd_sc_hd__nor3_2 _13800_ (.A(_08395_),
    .B(_08397_),
    .C(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__mux2i_2 _13801_ (.A0(net3719),
    .A1(_08357_),
    .S(_08348_),
    .Y(_08400_));
 sky130_fd_sc_hd__nand2_1 _13802_ (.A(_08205_),
    .B(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__o21ai_0 _13803_ (.A1(net3744),
    .A2(_08399_),
    .B1(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__a21oi_2 _13804_ (.A1(_08242_),
    .A2(_08359_),
    .B1(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__inv_2 _13805_ (.A(\cs_registers_i.pc_id_i[3] ),
    .Y(_08404_));
 sky130_fd_sc_hd__nand3_4 _13806_ (.A(net3833),
    .B(net337),
    .C(_08040_),
    .Y(_08405_));
 sky130_fd_sc_hd__nor2_4 _13807_ (.A(_08405_),
    .B(net3785),
    .Y(_08406_));
 sky130_fd_sc_hd__nand3_1 _13808_ (.A(net3897),
    .B(net3721),
    .C(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__o211ai_1 _13809_ (.A1(_08404_),
    .A2(net3721),
    .B1(_08407_),
    .C1(net3666),
    .Y(_08408_));
 sky130_fd_sc_hd__or3_1 _13810_ (.A(_08192_),
    .B(net3721),
    .C(net3716),
    .X(_08409_));
 sky130_fd_sc_hd__o211ai_1 _13811_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_08194_),
    .B1(_08408_),
    .C1(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__nor2_2 _13812_ (.A(_07857_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__a31oi_2 _13813_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(net3756),
    .A3(_07864_),
    .B1(_08411_),
    .Y(_08412_));
 sky130_fd_sc_hd__and2_4 _13814_ (.A(_08403_),
    .B(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__clkinv_2 _13815_ (.A(\cs_registers_i.pc_id_i[2] ),
    .Y(_08414_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1117 ();
 sky130_fd_sc_hd__nand3_1 _13818_ (.A(net3901),
    .B(net3723),
    .C(_08406_),
    .Y(_08417_));
 sky130_fd_sc_hd__o211ai_1 _13819_ (.A1(_08414_),
    .A2(net3723),
    .B1(_08417_),
    .C1(net3666),
    .Y(_08418_));
 sky130_fd_sc_hd__mux2i_1 _13820_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .S(net3933),
    .Y(_08419_));
 sky130_fd_sc_hd__mux2i_1 _13821_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(net3933),
    .Y(_08420_));
 sky130_fd_sc_hd__a221oi_1 _13822_ (.A1(net3793),
    .A2(_08419_),
    .B1(_08420_),
    .B2(net3791),
    .C1(net3896),
    .Y(_08421_));
 sky130_fd_sc_hd__mux2_1 _13823_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net3933),
    .X(_08422_));
 sky130_fd_sc_hd__a221o_1 _13824_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .A2(net3788),
    .B1(_08422_),
    .B2(net3915),
    .C1(_08160_),
    .X(_08423_));
 sky130_fd_sc_hd__o21ai_2 _13825_ (.A1(net350),
    .A2(_08421_),
    .B1(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__mux4_2 _13826_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S0(net3925),
    .S1(net3909),
    .X(_08425_));
 sky130_fd_sc_hd__mux4_2 _13827_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S0(net3925),
    .S1(net3909),
    .X(_08426_));
 sky130_fd_sc_hd__a22oi_2 _13828_ (.A1(_08126_),
    .A2(_08425_),
    .B1(_08426_),
    .B2(_08135_),
    .Y(_08427_));
 sky130_fd_sc_hd__mux4_2 _13829_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net3929),
    .S1(net3913),
    .X(_08428_));
 sky130_fd_sc_hd__mux4_2 _13830_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net3929),
    .S1(net3909),
    .X(_08429_));
 sky130_fd_sc_hd__mux4_2 _13831_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S0(net3925),
    .S1(net3909),
    .X(_08430_));
 sky130_fd_sc_hd__a22o_4 _13832_ (.A1(_08126_),
    .A2(_08429_),
    .B1(_08430_),
    .B2(net3796),
    .X(_08431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1116 ();
 sky130_fd_sc_hd__mux2i_1 _13834_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .S(net439),
    .Y(_08433_));
 sky130_fd_sc_hd__mux2i_1 _13835_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S(net439),
    .Y(_08434_));
 sky130_fd_sc_hd__o221ai_2 _13836_ (.A1(_08113_),
    .A2(_08433_),
    .B1(_08434_),
    .B2(_08119_),
    .C1(net3899),
    .Y(_08435_));
 sky130_fd_sc_hd__a211oi_4 _13837_ (.A1(_08111_),
    .A2(_08428_),
    .B1(_08431_),
    .C1(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__a21oi_4 _13838_ (.A1(_08427_),
    .A2(_08424_),
    .B1(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__or3_1 _13839_ (.A(_08192_),
    .B(net293),
    .C(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__o211ai_1 _13840_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(_08194_),
    .B1(_08418_),
    .C1(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand3_1 _13841_ (.A(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B(_07857_),
    .C(_07864_),
    .Y(_08440_));
 sky130_fd_sc_hd__o21ai_2 _13842_ (.A1(_08439_),
    .A2(_08316_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__nand2_8 _13843_ (.A(net300),
    .B(net3744),
    .Y(_08442_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1114 ();
 sky130_fd_sc_hd__nor3_1 _13846_ (.A(_07927_),
    .B(_07892_),
    .C(_08352_),
    .Y(_08445_));
 sky130_fd_sc_hd__a211oi_2 _13847_ (.A1(_07910_),
    .A2(_07908_),
    .B1(_08355_),
    .C1(net3947),
    .Y(_08446_));
 sky130_fd_sc_hd__o21ai_4 _13848_ (.A1(_08445_),
    .A2(_08446_),
    .B1(net3740),
    .Y(_08447_));
 sky130_fd_sc_hd__nand2_4 _13849_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(_08356_),
    .Y(_08448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1112 ();
 sky130_fd_sc_hd__mux4_2 _13852_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net3884),
    .S1(net3867),
    .X(_08451_));
 sky130_fd_sc_hd__nand2_1 _13853_ (.A(net3850),
    .B(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__mux4_2 _13854_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S0(net3884),
    .S1(net3867),
    .X(_08453_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(_07927_),
    .B(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__and3_4 _13856_ (.A(net3848),
    .B(_08452_),
    .C(_08454_),
    .X(_08455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1111 ();
 sky130_fd_sc_hd__mux2_1 _13858_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .S(net3850),
    .X(_08457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1109 ();
 sky130_fd_sc_hd__a22o_1 _13861_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .A2(net395),
    .B1(_08457_),
    .B2(net3867),
    .X(_08460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1106 ();
 sky130_fd_sc_hd__mux2i_1 _13865_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net3867),
    .Y(_08464_));
 sky130_fd_sc_hd__mux2i_1 _13866_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(net3867),
    .Y(_08465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1105 ();
 sky130_fd_sc_hd__o221ai_1 _13868_ (.A1(_07945_),
    .A2(_08464_),
    .B1(_08465_),
    .B2(_07951_),
    .C1(_07955_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21oi_1 _13869_ (.A1(_07935_),
    .A2(_08460_),
    .B1(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1102 ();
 sky130_fd_sc_hd__mux2i_1 _13873_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S(net3874),
    .Y(_08472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1101 ();
 sky130_fd_sc_hd__mux2i_1 _13875_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .S(net3874),
    .Y(_08474_));
 sky130_fd_sc_hd__a22oi_1 _13876_ (.A1(net3810),
    .A2(_08472_),
    .B1(_08474_),
    .B2(net3809),
    .Y(_08475_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1100 ();
 sky130_fd_sc_hd__mux2i_1 _13878_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .S(net3874),
    .Y(_08477_));
 sky130_fd_sc_hd__mux2i_1 _13879_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S(net3874),
    .Y(_08478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1099 ();
 sky130_fd_sc_hd__a22oi_1 _13881_ (.A1(net3804),
    .A2(_08477_),
    .B1(_08478_),
    .B2(net3803),
    .Y(_08480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1098 ();
 sky130_fd_sc_hd__mux4_2 _13883_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net3891),
    .S1(net3866),
    .X(_08482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1097 ();
 sky130_fd_sc_hd__mux4_2 _13885_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S0(net3891),
    .S1(net3866),
    .X(_08484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1096 ();
 sky130_fd_sc_hd__a22o_4 _13887_ (.A1(net3798),
    .A2(_08482_),
    .B1(_08484_),
    .B2(_07987_),
    .X(_08486_));
 sky130_fd_sc_hd__a31oi_4 _13888_ (.A1(net3751),
    .A2(_08475_),
    .A3(_08480_),
    .B1(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__o31ai_4 _13889_ (.A1(net3846),
    .A2(_08455_),
    .A3(_08468_),
    .B1(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nor2_2 _13890_ (.A(_08348_),
    .B(net3715),
    .Y(_08489_));
 sky130_fd_sc_hd__a41o_4 _13891_ (.A1(net3749),
    .A2(_08348_),
    .A3(_08447_),
    .A4(_08448_),
    .B1(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1095 ();
 sky130_fd_sc_hd__o22a_1 _13893_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .B2(net3787),
    .X(_08492_));
 sky130_fd_sc_hd__o221a_1 _13894_ (.A1(_08168_),
    .A2(_08437_),
    .B1(net3715),
    .B2(_08172_),
    .C1(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__nor2_1 _13895_ (.A(net3744),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__a21oi_2 _13896_ (.A1(_08205_),
    .A2(_08490_),
    .B1(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__o21ai_2 _13897_ (.A1(_08442_),
    .A2(_08490_),
    .B1(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__nor2_2 _13898_ (.A(_08496_),
    .B(_08441_),
    .Y(_08497_));
 sky130_fd_sc_hd__or3_4 _13899_ (.A(_08038_),
    .B(_07880_),
    .C(_08315_),
    .X(_08498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1094 ();
 sky130_fd_sc_hd__inv_12 _13901_ (.A(net3910),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_8 _13902_ (.A(_08188_),
    .B(_08075_),
    .Y(_08501_));
 sky130_fd_sc_hd__nor2_1 _13903_ (.A(_08500_),
    .B(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__mux2i_1 _13904_ (.A0(\cs_registers_i.pc_id_i[1] ),
    .A1(_08502_),
    .S(net293),
    .Y(_08503_));
 sky130_fd_sc_hd__mux2i_1 _13905_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .S(net3922),
    .Y(_08504_));
 sky130_fd_sc_hd__mux2i_1 _13906_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S(net3922),
    .Y(_08505_));
 sky130_fd_sc_hd__nor3_1 _13907_ (.A(_08109_),
    .B(_08504_),
    .C(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__mux2i_1 _13908_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .S(net3922),
    .Y(_08507_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1093 ();
 sky130_fd_sc_hd__mux2i_1 _13910_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S(net3922),
    .Y(_08509_));
 sky130_fd_sc_hd__nor3_1 _13911_ (.A(net3902),
    .B(_08507_),
    .C(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__mux4_2 _13912_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net3922),
    .S1(net3902),
    .X(_08511_));
 sky130_fd_sc_hd__mux4_2 _13913_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .S0(net3922),
    .S1(net3902),
    .X(_08512_));
 sky130_fd_sc_hd__mux2_1 _13914_ (.A0(_08511_),
    .A1(_08512_),
    .S(_08500_),
    .X(_08513_));
 sky130_fd_sc_hd__nor4_2 _13915_ (.A(_08287_),
    .B(_08506_),
    .C(_08510_),
    .D(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__mux2i_1 _13916_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .S(net3926),
    .Y(_08515_));
 sky130_fd_sc_hd__mux2i_1 _13917_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(net3926),
    .Y(_08516_));
 sky130_fd_sc_hd__a22oi_1 _13918_ (.A1(net3795),
    .A2(_08515_),
    .B1(_08516_),
    .B2(net412),
    .Y(_08517_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1092 ();
 sky130_fd_sc_hd__mux2i_1 _13920_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .S(net3926),
    .Y(_08519_));
 sky130_fd_sc_hd__mux2i_1 _13921_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S(net3926),
    .Y(_08520_));
 sky130_fd_sc_hd__a22oi_1 _13922_ (.A1(net478),
    .A2(_08519_),
    .B1(_08520_),
    .B2(net3778),
    .Y(_08521_));
 sky130_fd_sc_hd__nand2b_4 _13923_ (.A_N(net3899),
    .B(net3896),
    .Y(_08522_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1091 ();
 sky130_fd_sc_hd__a21oi_1 _13925_ (.A1(_08517_),
    .A2(_08521_),
    .B1(_08522_),
    .Y(_08524_));
 sky130_fd_sc_hd__mux2i_1 _13926_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .S(net3926),
    .Y(_08525_));
 sky130_fd_sc_hd__mux2i_1 _13927_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S(net3926),
    .Y(_08526_));
 sky130_fd_sc_hd__a22oi_1 _13928_ (.A1(net3795),
    .A2(_08525_),
    .B1(_08526_),
    .B2(net412),
    .Y(_08527_));
 sky130_fd_sc_hd__mux2i_1 _13929_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .S(net3926),
    .Y(_08528_));
 sky130_fd_sc_hd__mux2i_1 _13930_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S(net3926),
    .Y(_08529_));
 sky130_fd_sc_hd__a22oi_1 _13931_ (.A1(_08292_),
    .A2(_08528_),
    .B1(_08529_),
    .B2(net3778),
    .Y(_08530_));
 sky130_fd_sc_hd__nand2b_4 _13932_ (.A_N(net3896),
    .B(net3898),
    .Y(_08531_));
 sky130_fd_sc_hd__a21oi_1 _13933_ (.A1(_08527_),
    .A2(_08530_),
    .B1(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__mux2i_1 _13934_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .S(net3931),
    .Y(_08533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1090 ();
 sky130_fd_sc_hd__nand3b_1 _13936_ (.A_N(net3903),
    .B(net3931),
    .C(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .Y(_08535_));
 sky130_fd_sc_hd__o21ai_2 _13937_ (.A1(_08109_),
    .A2(_08533_),
    .B1(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__mux4_2 _13938_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S0(net3931),
    .S1(net3903),
    .X(_08537_));
 sky130_fd_sc_hd__or2_4 _13939_ (.A(net3896),
    .B(net349),
    .X(_08538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1089 ();
 sky130_fd_sc_hd__a21o_1 _13941_ (.A1(net3913),
    .A2(_08537_),
    .B1(_08538_),
    .X(_08540_));
 sky130_fd_sc_hd__a21oi_4 _13942_ (.A1(_08500_),
    .A2(_08536_),
    .B1(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__nor4_2 _13943_ (.A(_08514_),
    .B(_08524_),
    .C(_08532_),
    .D(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor3_2 _13944_ (.A(_08192_),
    .B(net293),
    .C(net3713),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_2 _13945_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .B(_08194_),
    .Y(_08544_));
 sky130_fd_sc_hd__a211oi_4 _13946_ (.A1(_08192_),
    .A2(_08503_),
    .B1(_08544_),
    .C1(_08543_),
    .Y(_08545_));
 sky130_fd_sc_hd__and3_4 _13947_ (.A(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .B(_07857_),
    .C(_07864_),
    .X(_08546_));
 sky130_fd_sc_hd__a21oi_2 _13948_ (.A1(_08498_),
    .A2(_08545_),
    .B1(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1088 ();
 sky130_fd_sc_hd__a211oi_1 _13950_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .A2(net296),
    .B1(net3849),
    .C1(net3893),
    .Y(_08549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1087 ();
 sky130_fd_sc_hd__mux2_1 _13952_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .S(net3854),
    .X(_08551_));
 sky130_fd_sc_hd__nand2_1 _13953_ (.A(net3879),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__mux4_2 _13954_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S0(net3879),
    .S1(net3854),
    .X(_08553_));
 sky130_fd_sc_hd__nor2_1 _13955_ (.A(_07935_),
    .B(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__a221oi_2 _13956_ (.A1(_08549_),
    .A2(_08552_),
    .B1(_08554_),
    .B2(_07955_),
    .C1(net3847),
    .Y(_08555_));
 sky130_fd_sc_hd__mux4_2 _13957_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S0(net404),
    .S1(net3854),
    .X(_08556_));
 sky130_fd_sc_hd__nor2_1 _13958_ (.A(net3893),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__mux4_2 _13959_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S0(net404),
    .S1(net3854),
    .X(_08558_));
 sky130_fd_sc_hd__nor3_1 _13960_ (.A(_07955_),
    .B(_07935_),
    .C(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__a21oi_1 _13961_ (.A1(net3849),
    .A2(_08557_),
    .B1(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__mux2i_1 _13962_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .S(net434),
    .Y(_08561_));
 sky130_fd_sc_hd__mux2i_2 _13963_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S(net434),
    .Y(_08562_));
 sky130_fd_sc_hd__a22oi_1 _13964_ (.A1(_07969_),
    .A2(_08561_),
    .B1(_08562_),
    .B2(_07962_),
    .Y(_08563_));
 sky130_fd_sc_hd__mux2i_1 _13965_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(net434),
    .Y(_08564_));
 sky130_fd_sc_hd__mux2i_1 _13966_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .S(net434),
    .Y(_08565_));
 sky130_fd_sc_hd__a22oi_2 _13967_ (.A1(_07983_),
    .A2(_08564_),
    .B1(_08565_),
    .B2(net312),
    .Y(_08566_));
 sky130_fd_sc_hd__and3_4 _13968_ (.A(_07960_),
    .B(_08563_),
    .C(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__mux2i_1 _13969_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(net3878),
    .Y(_08568_));
 sky130_fd_sc_hd__mux2i_1 _13970_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S(net3878),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2b_4 _13971_ (.A_N(net3884),
    .B(net3850),
    .Y(_08570_));
 sky130_fd_sc_hd__o22ai_1 _13972_ (.A1(_07951_),
    .A2(_08568_),
    .B1(_08569_),
    .B2(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__mux4_2 _13973_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S0(net3893),
    .S1(net3878),
    .X(_08572_));
 sky130_fd_sc_hd__a32o_1 _13974_ (.A1(net3847),
    .A2(net3849),
    .A3(_08571_),
    .B1(_08572_),
    .B2(net351),
    .X(_08573_));
 sky130_fd_sc_hd__a211oi_2 _13975_ (.A1(_08560_),
    .A2(_08555_),
    .B1(_08567_),
    .C1(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1084 ();
 sky130_fd_sc_hd__a21oi_4 _13979_ (.A1(_07908_),
    .A2(_07910_),
    .B1(net3754),
    .Y(_08578_));
 sky130_fd_sc_hd__mux2i_4 _13980_ (.A0(net3895),
    .A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .S(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__nand3_2 _13981_ (.A(_08348_),
    .B(net3740),
    .C(_07904_),
    .Y(_08580_));
 sky130_fd_sc_hd__o22a_4 _13982_ (.A1(_08348_),
    .A2(net3712),
    .B1(_08579_),
    .B2(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1081 ();
 sky130_fd_sc_hd__nand3_1 _13986_ (.A(net3933),
    .B(net293),
    .C(_08406_),
    .Y(_08585_));
 sky130_fd_sc_hd__mux2i_1 _13987_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(net3926),
    .Y(_08586_));
 sky130_fd_sc_hd__mux2i_1 _13988_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .S(net3926),
    .Y(_08587_));
 sky130_fd_sc_hd__a22o_1 _13989_ (.A1(_08147_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08292_),
    .X(_08588_));
 sky130_fd_sc_hd__mux2_1 _13990_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S(net3926),
    .X(_08589_));
 sky130_fd_sc_hd__mux2_1 _13991_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .S(net3926),
    .X(_08590_));
 sky130_fd_sc_hd__o22ai_1 _13992_ (.A1(_08266_),
    .A2(_08589_),
    .B1(_08590_),
    .B2(_08374_),
    .Y(_08591_));
 sky130_fd_sc_hd__o21ai_2 _13993_ (.A1(_08588_),
    .A2(_08591_),
    .B1(_08299_),
    .Y(_08592_));
 sky130_fd_sc_hd__mux2_1 _13994_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .S(net3926),
    .X(_08593_));
 sky130_fd_sc_hd__nand2b_1 _13995_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .B(net3926),
    .Y(_08594_));
 sky130_fd_sc_hd__o221ai_1 _13996_ (.A1(net3926),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .B1(_08593_),
    .B2(net3912),
    .C1(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__mux2_1 _13997_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .S(net3926),
    .X(_08596_));
 sky130_fd_sc_hd__mux2_1 _13998_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(net3926),
    .X(_08597_));
 sky130_fd_sc_hd__o211ai_1 _13999_ (.A1(net3912),
    .A2(_08596_),
    .B1(_08597_),
    .C1(net3903),
    .Y(_08598_));
 sky130_fd_sc_hd__a221oi_1 _14000_ (.A1(net263),
    .A2(_08596_),
    .B1(_08593_),
    .B2(net478),
    .C1(_08287_),
    .Y(_08599_));
 sky130_fd_sc_hd__o211ai_1 _14001_ (.A1(net3903),
    .A2(_08595_),
    .B1(_08598_),
    .C1(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__mux2i_1 _14002_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(net3927),
    .Y(_08601_));
 sky130_fd_sc_hd__mux2i_1 _14003_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .S(net3927),
    .Y(_08602_));
 sky130_fd_sc_hd__o22ai_1 _14004_ (.A1(_08261_),
    .A2(_08601_),
    .B1(_08602_),
    .B2(_08374_),
    .Y(_08603_));
 sky130_fd_sc_hd__nor3b_4 _14005_ (.A(net3902),
    .B(net3908),
    .C_N(net3927),
    .Y(_08604_));
 sky130_fd_sc_hd__mux2i_1 _14006_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net3927),
    .Y(_08605_));
 sky130_fd_sc_hd__o2bb2ai_1 _14007_ (.A1_N(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .A2_N(_08604_),
    .B1(_08605_),
    .B2(_08266_),
    .Y(_08606_));
 sky130_fd_sc_hd__or3_4 _14008_ (.A(_08538_),
    .B(_08603_),
    .C(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__mux2_1 _14009_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .S(net3926),
    .X(_08608_));
 sky130_fd_sc_hd__nand2b_1 _14010_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .B(net3926),
    .Y(_08609_));
 sky130_fd_sc_hd__o221ai_1 _14011_ (.A1(net3926),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .B1(_08608_),
    .B2(net3912),
    .C1(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__mux2_1 _14012_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .S(net3926),
    .X(_08611_));
 sky130_fd_sc_hd__mux2_1 _14013_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(net3926),
    .X(_08612_));
 sky130_fd_sc_hd__o211ai_1 _14014_ (.A1(net3912),
    .A2(_08611_),
    .B1(_08612_),
    .C1(net3903),
    .Y(_08613_));
 sky130_fd_sc_hd__a221oi_1 _14015_ (.A1(net263),
    .A2(_08611_),
    .B1(_08608_),
    .B2(net259),
    .C1(_08531_),
    .Y(_08614_));
 sky130_fd_sc_hd__o211ai_1 _14016_ (.A1(net3903),
    .A2(_08610_),
    .B1(_08613_),
    .C1(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__nand4_1 _14017_ (.A(_08592_),
    .B(_08600_),
    .C(_08607_),
    .D(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__inv_1 _14018_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .Y(_08617_));
 sky130_fd_sc_hd__mux2_1 _14019_ (.A0(net3709),
    .A1(_08617_),
    .S(net293),
    .X(_08618_));
 sky130_fd_sc_hd__nand2b_4 _14020_ (.A_N(_08191_),
    .B(_08194_),
    .Y(_08619_));
 sky130_fd_sc_hd__mux2_8 _14021_ (.A0(_08585_),
    .A1(_08618_),
    .S(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_2 _14022_ (.A(_08581_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand2_2 _14023_ (.A(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .B(_07864_),
    .Y(_08622_));
 sky130_fd_sc_hd__nor3_4 _14024_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .C(_07864_),
    .Y(_08623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1079 ();
 sky130_fd_sc_hd__o22ai_1 _14027_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .B2(net3787),
    .Y(_08626_));
 sky130_fd_sc_hd__a221oi_4 _14028_ (.A1(_08623_),
    .A2(net3712),
    .B1(net3710),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .C1(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__a21oi_2 _14029_ (.A1(_08622_),
    .A2(_08627_),
    .B1(_08498_),
    .Y(_08628_));
 sky130_fd_sc_hd__o22ai_2 _14030_ (.A1(_08348_),
    .A2(net3712),
    .B1(_08579_),
    .B2(_08580_),
    .Y(_08629_));
 sky130_fd_sc_hd__nor2_1 _14031_ (.A(_08095_),
    .B(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__a211oi_2 _14032_ (.A1(net3744),
    .A2(_08621_),
    .B1(_08628_),
    .C1(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_4 _14033_ (.A(_07887_),
    .B(_07910_),
    .Y(_08632_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1077 ();
 sky130_fd_sc_hd__nor2b_1 _14036_ (.A(_08355_),
    .B_N(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Y(_08635_));
 sky130_fd_sc_hd__mux2i_1 _14037_ (.A0(net3858),
    .A1(_08635_),
    .S(_08578_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _14038_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .B(_08356_),
    .Y(_08637_));
 sky130_fd_sc_hd__o21ai_2 _14039_ (.A1(_08632_),
    .A2(_08636_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__mux4_2 _14040_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S0(net3893),
    .S1(net3875),
    .X(_08639_));
 sky130_fd_sc_hd__nand2_2 _14041_ (.A(net3854),
    .B(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__mux4_2 _14042_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S0(net3893),
    .S1(net3875),
    .X(_08641_));
 sky130_fd_sc_hd__nand2_2 _14043_ (.A(_07927_),
    .B(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__nand3_4 _14044_ (.A(net3848),
    .B(_08640_),
    .C(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__mux2_1 _14045_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .S(net3850),
    .X(_08644_));
 sky130_fd_sc_hd__a22o_1 _14046_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .A2(net3816),
    .B1(_08644_),
    .B2(net303),
    .X(_08645_));
 sky130_fd_sc_hd__mux2i_1 _14047_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net3867),
    .Y(_08646_));
 sky130_fd_sc_hd__mux2i_1 _14048_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(net3867),
    .Y(_08647_));
 sky130_fd_sc_hd__o22ai_1 _14049_ (.A1(_07945_),
    .A2(_08646_),
    .B1(_08647_),
    .B2(_07951_),
    .Y(_08648_));
 sky130_fd_sc_hd__a211o_4 _14050_ (.A1(_07935_),
    .A2(_08645_),
    .B1(_08648_),
    .C1(net3849),
    .X(_08649_));
 sky130_fd_sc_hd__nand2b_4 _14051_ (.A_N(net3849),
    .B(net3847),
    .Y(_08650_));
 sky130_fd_sc_hd__mux2_4 _14052_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S(net434),
    .X(_08651_));
 sky130_fd_sc_hd__mux2_1 _14053_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .S(net434),
    .X(_08652_));
 sky130_fd_sc_hd__o22ai_2 _14054_ (.A1(net361),
    .A2(_08651_),
    .B1(_08652_),
    .B2(_08570_),
    .Y(_08653_));
 sky130_fd_sc_hd__mux2i_1 _14055_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .S(net434),
    .Y(_08654_));
 sky130_fd_sc_hd__mux2i_1 _14056_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(net434),
    .Y(_08655_));
 sky130_fd_sc_hd__a22o_4 _14057_ (.A1(net312),
    .A2(_08654_),
    .B1(_08655_),
    .B2(net3802),
    .X(_08656_));
 sky130_fd_sc_hd__mux4_2 _14058_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S0(net3888),
    .S1(net434),
    .X(_08657_));
 sky130_fd_sc_hd__mux4_2 _14059_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net3888),
    .S1(net434),
    .X(_08658_));
 sky130_fd_sc_hd__a22oi_2 _14060_ (.A1(net351),
    .A2(_08657_),
    .B1(_08658_),
    .B2(net3798),
    .Y(_08659_));
 sky130_fd_sc_hd__o31ai_4 _14061_ (.A1(_08650_),
    .A2(_08653_),
    .A3(_08656_),
    .B1(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__a31oi_4 _14062_ (.A1(_08649_),
    .A2(_08643_),
    .A3(_07958_),
    .B1(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__nor2_1 _14063_ (.A(_08348_),
    .B(net342),
    .Y(_08662_));
 sky130_fd_sc_hd__a21o_4 _14064_ (.A1(_08348_),
    .A2(_08638_),
    .B1(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__a211oi_2 _14065_ (.A1(_08348_),
    .A2(_08638_),
    .B1(_08662_),
    .C1(_08095_),
    .Y(_08664_));
 sky130_fd_sc_hd__o22ai_1 _14066_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .B2(net3787),
    .Y(_08665_));
 sky130_fd_sc_hd__a21oi_1 _14067_ (.A1(_08623_),
    .A2(net342),
    .B1(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__o21a_1 _14068_ (.A1(_08168_),
    .A2(net3713),
    .B1(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__nor2_1 _14069_ (.A(net3748),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__a211oi_4 _14070_ (.A1(_08242_),
    .A2(_08663_),
    .B1(_08664_),
    .C1(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__maj3_2 _14071_ (.A(_08547_),
    .B(_08669_),
    .C(_08631_),
    .X(_08670_));
 sky130_fd_sc_hd__nand2_2 _14072_ (.A(_08441_),
    .B(_08496_),
    .Y(_08671_));
 sky130_fd_sc_hd__o221a_4 _14073_ (.A1(_08403_),
    .A2(_08412_),
    .B1(_08497_),
    .B2(_08670_),
    .C1(_08671_),
    .X(_08672_));
 sky130_fd_sc_hd__mux2i_1 _14074_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .S(net3924),
    .Y(_08673_));
 sky130_fd_sc_hd__mux2i_1 _14075_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(net3924),
    .Y(_08674_));
 sky130_fd_sc_hd__a22oi_1 _14076_ (.A1(net3776),
    .A2(_08673_),
    .B1(_08674_),
    .B2(_08147_),
    .Y(_08675_));
 sky130_fd_sc_hd__mux2i_1 _14077_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .S(net3924),
    .Y(_08676_));
 sky130_fd_sc_hd__mux2i_1 _14078_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S(net3924),
    .Y(_08677_));
 sky130_fd_sc_hd__a22oi_1 _14079_ (.A1(net3795),
    .A2(_08676_),
    .B1(_08677_),
    .B2(net3778),
    .Y(_08678_));
 sky130_fd_sc_hd__nand3_1 _14080_ (.A(net3784),
    .B(_08675_),
    .C(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__mux2i_1 _14081_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(net3923),
    .Y(_08680_));
 sky130_fd_sc_hd__mux2i_1 _14082_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net3923),
    .Y(_08681_));
 sky130_fd_sc_hd__o22ai_1 _14083_ (.A1(_08261_),
    .A2(_08680_),
    .B1(_08681_),
    .B2(_08266_),
    .Y(_08682_));
 sky130_fd_sc_hd__mux2i_1 _14084_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .S(net3923),
    .Y(_08683_));
 sky130_fd_sc_hd__a21oi_1 _14085_ (.A1(net3923),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B1(net3902),
    .Y(_08684_));
 sky130_fd_sc_hd__a211oi_1 _14086_ (.A1(net3902),
    .A2(_08683_),
    .B1(_08684_),
    .C1(net3910),
    .Y(_08685_));
 sky130_fd_sc_hd__o21ai_2 _14087_ (.A1(_08682_),
    .A2(_08685_),
    .B1(net3781),
    .Y(_08686_));
 sky130_fd_sc_hd__mux2i_1 _14088_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .S(net3924),
    .Y(_08687_));
 sky130_fd_sc_hd__mux2i_1 _14089_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .S(net3924),
    .Y(_08688_));
 sky130_fd_sc_hd__a22oi_1 _14090_ (.A1(net3776),
    .A2(_08687_),
    .B1(_08688_),
    .B2(net3795),
    .Y(_08689_));
 sky130_fd_sc_hd__mux2i_1 _14091_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S(net3924),
    .Y(_08690_));
 sky130_fd_sc_hd__mux2i_1 _14092_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S(net3924),
    .Y(_08691_));
 sky130_fd_sc_hd__a22oi_1 _14093_ (.A1(_08147_),
    .A2(_08690_),
    .B1(_08691_),
    .B2(net3778),
    .Y(_08692_));
 sky130_fd_sc_hd__nand3_1 _14094_ (.A(net3774),
    .B(_08689_),
    .C(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__and2_4 _14095_ (.A(net3896),
    .B(net3898),
    .X(_08694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1076 ();
 sky130_fd_sc_hd__mux2i_1 _14097_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S(net3924),
    .Y(_08696_));
 sky130_fd_sc_hd__mux2i_1 _14098_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .S(net3924),
    .Y(_08697_));
 sky130_fd_sc_hd__a22oi_1 _14099_ (.A1(net3778),
    .A2(_08696_),
    .B1(_08697_),
    .B2(net3795),
    .Y(_08698_));
 sky130_fd_sc_hd__mux2i_1 _14100_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .S(net3924),
    .Y(_08699_));
 sky130_fd_sc_hd__mux2i_1 _14101_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S(net3924),
    .Y(_08700_));
 sky130_fd_sc_hd__a22oi_1 _14102_ (.A1(net3776),
    .A2(_08699_),
    .B1(_08700_),
    .B2(_08147_),
    .Y(_08701_));
 sky130_fd_sc_hd__nand3_1 _14103_ (.A(_08694_),
    .B(_08698_),
    .C(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__and4_4 _14104_ (.A(_08693_),
    .B(_08686_),
    .C(_08679_),
    .D(_08702_),
    .X(_08703_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1075 ();
 sky130_fd_sc_hd__nand2b_2 _14106_ (.A_N(net3721),
    .B(_08703_),
    .Y(_08705_));
 sky130_fd_sc_hd__inv_1 _14107_ (.A(\cs_registers_i.pc_id_i[4] ),
    .Y(_08706_));
 sky130_fd_sc_hd__nand3_1 _14108_ (.A(net3896),
    .B(net3721),
    .C(_08406_),
    .Y(_08707_));
 sky130_fd_sc_hd__o211ai_1 _14109_ (.A1(_08706_),
    .A2(net3721),
    .B1(_08707_),
    .C1(net3666),
    .Y(_08708_));
 sky130_fd_sc_hd__o221ai_4 _14110_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(_08194_),
    .B1(net270),
    .B2(_08705_),
    .C1(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__nor2_1 _14111_ (.A(net3756),
    .B(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__a31oi_2 _14112_ (.A1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A2(net3756),
    .A3(_07864_),
    .B1(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__mux4_2 _14113_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S0(net3889),
    .S1(net3865),
    .X(_08712_));
 sky130_fd_sc_hd__nand2_1 _14114_ (.A(net3855),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__mux4_2 _14115_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S0(net3889),
    .S1(net3865),
    .X(_08714_));
 sky130_fd_sc_hd__nand2_1 _14116_ (.A(_07927_),
    .B(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__and3_4 _14117_ (.A(net3848),
    .B(_08713_),
    .C(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__mux2_1 _14118_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .S(net3855),
    .X(_08717_));
 sky130_fd_sc_hd__a22o_1 _14119_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .A2(net296),
    .B1(_08717_),
    .B2(net3875),
    .X(_08718_));
 sky130_fd_sc_hd__mux2i_1 _14120_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net3875),
    .Y(_08719_));
 sky130_fd_sc_hd__mux2i_1 _14121_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(net3875),
    .Y(_08720_));
 sky130_fd_sc_hd__o221ai_1 _14122_ (.A1(net363),
    .A2(_08719_),
    .B1(_08720_),
    .B2(net426),
    .C1(_07955_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21oi_1 _14123_ (.A1(_07935_),
    .A2(_08718_),
    .B1(_08721_),
    .Y(_08722_));
 sky130_fd_sc_hd__mux2i_1 _14124_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S(net3865),
    .Y(_08723_));
 sky130_fd_sc_hd__mux2i_1 _14125_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .S(net3865),
    .Y(_08724_));
 sky130_fd_sc_hd__a22oi_2 _14126_ (.A1(net3811),
    .A2(_08723_),
    .B1(_08724_),
    .B2(net3808),
    .Y(_08725_));
 sky130_fd_sc_hd__mux2i_1 _14127_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .S(net3865),
    .Y(_08726_));
 sky130_fd_sc_hd__mux2i_1 _14128_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S(net3865),
    .Y(_08727_));
 sky130_fd_sc_hd__a22oi_2 _14129_ (.A1(net312),
    .A2(_08726_),
    .B1(_08727_),
    .B2(net3802),
    .Y(_08728_));
 sky130_fd_sc_hd__mux4_2 _14130_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S0(net3888),
    .S1(net3865),
    .X(_08729_));
 sky130_fd_sc_hd__mux4_2 _14131_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S0(net3890),
    .S1(net3865),
    .X(_08730_));
 sky130_fd_sc_hd__a22o_1 _14132_ (.A1(net3798),
    .A2(_08729_),
    .B1(_08730_),
    .B2(net275),
    .X(_08731_));
 sky130_fd_sc_hd__a31oi_4 _14133_ (.A1(net3752),
    .A2(_08725_),
    .A3(_08728_),
    .B1(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__o31ai_2 _14134_ (.A1(net3844),
    .A2(_08716_),
    .A3(_08722_),
    .B1(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1074 ();
 sky130_fd_sc_hd__nor2_2 _14136_ (.A(_08632_),
    .B(_08578_),
    .Y(_08735_));
 sky130_fd_sc_hd__a22o_4 _14137_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_08356_),
    .B1(_08735_),
    .B2(net3845),
    .X(_08736_));
 sky130_fd_sc_hd__mux2_8 _14138_ (.A0(net3707),
    .A1(_08736_),
    .S(_08348_),
    .X(_08737_));
 sky130_fd_sc_hd__nor2_1 _14139_ (.A(_08172_),
    .B(net3707),
    .Y(_08738_));
 sky130_fd_sc_hd__o22ai_1 _14140_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .B2(net3787),
    .Y(_08739_));
 sky130_fd_sc_hd__a211oi_2 _14141_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_08703_),
    .B1(_08738_),
    .C1(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__o22ai_1 _14142_ (.A1(net299),
    .A2(_08737_),
    .B1(_08740_),
    .B2(net3748),
    .Y(_08741_));
 sky130_fd_sc_hd__a21oi_2 _14143_ (.A1(_08242_),
    .A2(_08737_),
    .B1(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__and2_0 _14144_ (.A(_08711_),
    .B(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__or2_0 _14145_ (.A(_08711_),
    .B(_08742_),
    .X(_08744_));
 sky130_fd_sc_hd__o31ai_4 _14146_ (.A1(_08413_),
    .A2(_08672_),
    .A3(_08743_),
    .B1(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__nand2_1 _14147_ (.A(net3756),
    .B(_07866_),
    .Y(_08746_));
 sky130_fd_sc_hd__o21ai_0 _14148_ (.A1(_08204_),
    .A2(_08316_),
    .B1(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1073 ();
 sky130_fd_sc_hd__mux2i_1 _14150_ (.A0(_08205_),
    .A1(net289),
    .S(_08000_),
    .Y(_08749_));
 sky130_fd_sc_hd__o21ai_0 _14151_ (.A1(net3748),
    .A2(_08178_),
    .B1(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__nand3_1 _14152_ (.A(net485),
    .B(_08319_),
    .C(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__a21oi_1 _14153_ (.A1(net485),
    .A2(_08319_),
    .B1(_08750_),
    .Y(_08752_));
 sky130_fd_sc_hd__a21oi_2 _14154_ (.A1(_08747_),
    .A2(_08751_),
    .B1(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__a31oi_4 _14155_ (.A1(_08210_),
    .A2(_08321_),
    .A3(_08745_),
    .B1(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__mux4_2 _14156_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net322),
    .S1(net303),
    .X(_08755_));
 sky130_fd_sc_hd__nand2_1 _14157_ (.A(net294),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__mux4_2 _14158_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S0(net322),
    .S1(net303),
    .X(_08757_));
 sky130_fd_sc_hd__nand2_1 _14159_ (.A(net3817),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__and3_4 _14160_ (.A(net3848),
    .B(_08756_),
    .C(_08758_),
    .X(_08759_));
 sky130_fd_sc_hd__mux2_1 _14161_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .S(net295),
    .X(_08760_));
 sky130_fd_sc_hd__a22o_4 _14162_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .A2(net3815),
    .B1(_08760_),
    .B2(net262),
    .X(_08761_));
 sky130_fd_sc_hd__mux2i_1 _14163_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net303),
    .Y(_08762_));
 sky130_fd_sc_hd__mux2i_1 _14164_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(net303),
    .Y(_08763_));
 sky130_fd_sc_hd__o22ai_2 _14165_ (.A1(net3814),
    .A2(_08762_),
    .B1(_08763_),
    .B2(net430),
    .Y(_08764_));
 sky130_fd_sc_hd__a211oi_4 _14166_ (.A1(_07935_),
    .A2(_08761_),
    .B1(_08764_),
    .C1(net3848),
    .Y(_08765_));
 sky130_fd_sc_hd__mux2i_1 _14167_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(net3876),
    .Y(_08766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1072 ();
 sky130_fd_sc_hd__mux2i_1 _14169_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .S(net3876),
    .Y(_08768_));
 sky130_fd_sc_hd__a22oi_1 _14170_ (.A1(net3810),
    .A2(_08766_),
    .B1(_08768_),
    .B2(net3809),
    .Y(_08769_));
 sky130_fd_sc_hd__mux2i_1 _14171_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .S(net3876),
    .Y(_08770_));
 sky130_fd_sc_hd__mux2i_1 _14172_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S(net3876),
    .Y(_08771_));
 sky130_fd_sc_hd__a22oi_1 _14173_ (.A1(net3804),
    .A2(_08770_),
    .B1(_08771_),
    .B2(net3803),
    .Y(_08772_));
 sky130_fd_sc_hd__mux4_2 _14174_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S0(net3884),
    .S1(net3876),
    .X(_08773_));
 sky130_fd_sc_hd__mux4_2 _14175_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net322),
    .S1(net3876),
    .X(_08774_));
 sky130_fd_sc_hd__a22o_4 _14176_ (.A1(net279),
    .A2(_08773_),
    .B1(_08774_),
    .B2(net3798),
    .X(_08775_));
 sky130_fd_sc_hd__a31oi_4 _14177_ (.A1(net3751),
    .A2(_08769_),
    .A3(_08772_),
    .B1(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__o31ai_4 _14178_ (.A1(_08759_),
    .A2(net3846),
    .A3(_08765_),
    .B1(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1071 ();
 sky130_fd_sc_hd__a22o_4 _14180_ (.A1(net3841),
    .A2(net3667),
    .B1(_08777_),
    .B2(net3728),
    .X(_08779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1070 ();
 sky130_fd_sc_hd__mux2i_1 _14182_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .S(net3934),
    .Y(_08781_));
 sky130_fd_sc_hd__mux2i_1 _14183_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(net3934),
    .Y(_08782_));
 sky130_fd_sc_hd__a221oi_2 _14184_ (.A1(net3793),
    .A2(_08781_),
    .B1(_08782_),
    .B2(net3791),
    .C1(net3896),
    .Y(_08783_));
 sky130_fd_sc_hd__mux2_1 _14185_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net3934),
    .X(_08784_));
 sky130_fd_sc_hd__a221o_1 _14186_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .A2(net3788),
    .B1(_08784_),
    .B2(net3915),
    .C1(_08160_),
    .X(_08785_));
 sky130_fd_sc_hd__o21ai_4 _14187_ (.A1(net350),
    .A2(_08783_),
    .B1(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__mux4_2 _14188_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S0(net3931),
    .S1(net3913),
    .X(_08787_));
 sky130_fd_sc_hd__mux4_2 _14189_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S0(net3931),
    .S1(net3913),
    .X(_08788_));
 sky130_fd_sc_hd__a22oi_2 _14190_ (.A1(_08126_),
    .A2(_08787_),
    .B1(_08788_),
    .B2(_08135_),
    .Y(_08789_));
 sky130_fd_sc_hd__mux4_2 _14191_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net309),
    .S1(net3916),
    .X(_08790_));
 sky130_fd_sc_hd__mux2i_1 _14192_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .S(net267),
    .Y(_08791_));
 sky130_fd_sc_hd__mux2i_1 _14193_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S(net267),
    .Y(_08792_));
 sky130_fd_sc_hd__o221ai_1 _14194_ (.A1(_08113_),
    .A2(_08791_),
    .B1(_08792_),
    .B2(_08119_),
    .C1(net3899),
    .Y(_08793_));
 sky130_fd_sc_hd__a21oi_2 _14195_ (.A1(_08126_),
    .A2(_08790_),
    .B1(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__mux4_2 _14196_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net439),
    .S1(net3916),
    .X(_08795_));
 sky130_fd_sc_hd__mux4_2 _14197_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S0(net3931),
    .S1(net3913),
    .X(_08796_));
 sky130_fd_sc_hd__a22oi_2 _14198_ (.A1(_08111_),
    .A2(_08795_),
    .B1(_08796_),
    .B2(_08135_),
    .Y(_08797_));
 sky130_fd_sc_hd__a22o_4 _14199_ (.A1(_08786_),
    .A2(_08789_),
    .B1(_08794_),
    .B2(_08797_),
    .X(_08798_));
 sky130_fd_sc_hd__o22ai_1 _14200_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .B2(net3787),
    .Y(_08799_));
 sky130_fd_sc_hd__nor2_1 _14201_ (.A(_08172_),
    .B(_08777_),
    .Y(_08800_));
 sky130_fd_sc_hd__a211oi_1 _14202_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net402),
    .B1(_08799_),
    .C1(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1069 ();
 sky130_fd_sc_hd__o22ai_2 _14204_ (.A1(net3747),
    .A2(_08801_),
    .B1(_08779_),
    .B2(net3626),
    .Y(_08803_));
 sky130_fd_sc_hd__a21oi_4 _14205_ (.A1(net3624),
    .A2(_08779_),
    .B1(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1067 ();
 sky130_fd_sc_hd__nor2_1 _14208_ (.A(net3721),
    .B(_08798_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21oi_1 _14209_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net3721),
    .B1(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_2 _14210_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(net3665),
    .Y(_08809_));
 sky130_fd_sc_hd__o21ai_4 _14211_ (.A1(net3666),
    .A2(_08808_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__and3_1 _14212_ (.A(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B(net3755),
    .C(_07864_),
    .X(_08811_));
 sky130_fd_sc_hd__a21oi_2 _14213_ (.A1(net3745),
    .A2(_08810_),
    .B1(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__xor2_2 _14214_ (.A(_08804_),
    .B(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__xnor2_4 _14215_ (.A(net3541),
    .B(_08813_),
    .Y(net178));
 sky130_fd_sc_hd__maj3_1 _14216_ (.A(net280),
    .B(_08319_),
    .C(net3553),
    .X(_08814_));
 sky130_fd_sc_hd__xnor2_2 _14217_ (.A(_08210_),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__inv_1 _14218_ (.A(net3529),
    .Y(net177));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1065 ();
 sky130_fd_sc_hd__nand2_2 _14221_ (.A(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B(_07864_),
    .Y(_08818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1064 ();
 sky130_fd_sc_hd__nor2b_4 _14223_ (.A(net3844),
    .B_N(net3849),
    .Y(_08820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1063 ();
 sky130_fd_sc_hd__mux4_2 _14225_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S0(net3888),
    .S1(net3864),
    .X(_08822_));
 sky130_fd_sc_hd__mux4_2 _14226_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S0(net3888),
    .S1(net3864),
    .X(_08823_));
 sky130_fd_sc_hd__mux2i_1 _14227_ (.A0(_08822_),
    .A1(_08823_),
    .S(_07927_),
    .Y(_08824_));
 sky130_fd_sc_hd__mux2i_1 _14228_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S(net359),
    .Y(_08825_));
 sky130_fd_sc_hd__mux2i_1 _14229_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .S(net359),
    .Y(_08826_));
 sky130_fd_sc_hd__a221oi_1 _14230_ (.A1(_07983_),
    .A2(_08825_),
    .B1(_08826_),
    .B2(_07969_),
    .C1(net3844),
    .Y(_08827_));
 sky130_fd_sc_hd__mux2_1 _14231_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net405),
    .X(_08828_));
 sky130_fd_sc_hd__nor2b_4 _14232_ (.A(net341),
    .B_N(net359),
    .Y(_08829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1062 ();
 sky130_fd_sc_hd__a221o_1 _14234_ (.A1(net3892),
    .A2(_08828_),
    .B1(_08829_),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .C1(net3854),
    .X(_08831_));
 sky130_fd_sc_hd__a21oi_2 _14235_ (.A1(_08827_),
    .A2(_08831_),
    .B1(net3848),
    .Y(_08832_));
 sky130_fd_sc_hd__mux4_2 _14236_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .S0(net3864),
    .S1(net3852),
    .X(_08833_));
 sky130_fd_sc_hd__nor2b_2 _14237_ (.A(net3888),
    .B_N(net3844),
    .Y(_08834_));
 sky130_fd_sc_hd__mux4_2 _14238_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S0(net359),
    .S1(net3852),
    .X(_08835_));
 sky130_fd_sc_hd__and3_1 _14239_ (.A(net3844),
    .B(net3888),
    .C(_08835_),
    .X(_08836_));
 sky130_fd_sc_hd__a21oi_2 _14240_ (.A1(_08833_),
    .A2(_08834_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1061 ();
 sky130_fd_sc_hd__nand2_8 _14242_ (.A(net3844),
    .B(net3848),
    .Y(_08839_));
 sky130_fd_sc_hd__mux4_2 _14243_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S0(net3882),
    .S1(net3860),
    .X(_08840_));
 sky130_fd_sc_hd__mux4_2 _14244_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net3882),
    .S1(net3860),
    .X(_08841_));
 sky130_fd_sc_hd__nand2b_1 _14245_ (.A_N(_08841_),
    .B(_07993_),
    .Y(_08842_));
 sky130_fd_sc_hd__o31ai_2 _14246_ (.A1(net3853),
    .A2(_08839_),
    .A3(_08840_),
    .B1(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__a221oi_4 _14247_ (.A1(net407),
    .A2(_08824_),
    .B1(_08837_),
    .B2(_08832_),
    .C1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__a22o_4 _14248_ (.A1(net3839),
    .A2(_07912_),
    .B1(net3706),
    .B2(_07888_),
    .X(_08845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1060 ();
 sky130_fd_sc_hd__mux2_1 _14250_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net346),
    .X(_08847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1059 ();
 sky130_fd_sc_hd__a221oi_2 _14252_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .A2(net319),
    .B1(_08847_),
    .B2(net3910),
    .C1(net3905),
    .Y(_08849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1058 ();
 sky130_fd_sc_hd__mux4_2 _14254_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net3925),
    .S1(net3908),
    .X(_08851_));
 sky130_fd_sc_hd__o21ai_0 _14255_ (.A1(_08109_),
    .A2(_08851_),
    .B1(_08279_),
    .Y(_08852_));
 sky130_fd_sc_hd__mux4_2 _14256_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S0(net396),
    .S1(net3906),
    .X(_08853_));
 sky130_fd_sc_hd__and3b_4 _14257_ (.A_N(net283),
    .B(net3898),
    .C(net3896),
    .X(_08854_));
 sky130_fd_sc_hd__and3_4 _14258_ (.A(net3896),
    .B(net3898),
    .C(net283),
    .X(_08855_));
 sky130_fd_sc_hd__mux4_2 _14259_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net396),
    .S1(net3906),
    .X(_08856_));
 sky130_fd_sc_hd__a22oi_1 _14260_ (.A1(_08853_),
    .A2(_08854_),
    .B1(_08855_),
    .B2(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__o21ai_0 _14261_ (.A1(_08849_),
    .A2(_08852_),
    .B1(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1056 ();
 sky130_fd_sc_hd__mux2i_1 _14264_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S(net3923),
    .Y(_08861_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1055 ();
 sky130_fd_sc_hd__mux2i_1 _14266_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .S(net3923),
    .Y(_08863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1054 ();
 sky130_fd_sc_hd__a22oi_1 _14268_ (.A1(net370),
    .A2(_08861_),
    .B1(_08863_),
    .B2(net263),
    .Y(_08865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1053 ();
 sky130_fd_sc_hd__mux2i_1 _14270_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .S(net3923),
    .Y(_08867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1051 ();
 sky130_fd_sc_hd__mux2i_1 _14273_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S(net3923),
    .Y(_08870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1050 ();
 sky130_fd_sc_hd__a22oi_1 _14275_ (.A1(net260),
    .A2(_08867_),
    .B1(_08870_),
    .B2(_08147_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand3_1 _14276_ (.A(net3772),
    .B(_08865_),
    .C(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__mux2i_1 _14277_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .S(net3923),
    .Y(_08874_));
 sky130_fd_sc_hd__mux2i_1 _14278_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .S(net3923),
    .Y(_08875_));
 sky130_fd_sc_hd__a22oi_1 _14279_ (.A1(net260),
    .A2(_08874_),
    .B1(_08875_),
    .B2(net264),
    .Y(_08876_));
 sky130_fd_sc_hd__mux2i_1 _14280_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S(net3923),
    .Y(_08877_));
 sky130_fd_sc_hd__mux2i_1 _14281_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(net3923),
    .Y(_08878_));
 sky130_fd_sc_hd__a22oi_1 _14282_ (.A1(net370),
    .A2(_08877_),
    .B1(_08878_),
    .B2(_08147_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand3_1 _14283_ (.A(_08258_),
    .B(_08876_),
    .C(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__and3b_4 _14284_ (.A_N(_08858_),
    .B(_08873_),
    .C(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__nor2_1 _14285_ (.A(_08172_),
    .B(net340),
    .Y(_08882_));
 sky130_fd_sc_hd__o22ai_1 _14286_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .B2(_08171_),
    .Y(_08883_));
 sky130_fd_sc_hd__a211oi_2 _14287_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_08881_),
    .B1(_08882_),
    .C1(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__o21ai_0 _14288_ (.A1(net3626),
    .A2(_08845_),
    .B1(net473),
    .Y(_08885_));
 sky130_fd_sc_hd__xor2_1 _14289_ (.A(_08818_),
    .B(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1049 ();
 sky130_fd_sc_hd__inv_1 _14291_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .Y(_08888_));
 sky130_fd_sc_hd__mux2i_1 _14292_ (.A0(_08881_),
    .A1(_08888_),
    .S(net3720),
    .Y(_08889_));
 sky130_fd_sc_hd__a22o_4 _14293_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(_08202_),
    .B1(_08889_),
    .B2(net483),
    .X(_08890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1048 ();
 sky130_fd_sc_hd__xnor2_1 _14295_ (.A(_08845_),
    .B(net3617),
    .Y(_08892_));
 sky130_fd_sc_hd__xnor2_1 _14296_ (.A(_08205_),
    .B(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__nor2_1 _14297_ (.A(_07857_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__a21oi_2 _14298_ (.A1(_07857_),
    .A2(_08886_),
    .B1(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__nand2_2 _14299_ (.A(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .B(_07864_),
    .Y(_08896_));
 sky130_fd_sc_hd__mux2i_1 _14300_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .S(net3879),
    .Y(_08897_));
 sky130_fd_sc_hd__mux2i_1 _14301_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S(net3879),
    .Y(_08898_));
 sky130_fd_sc_hd__a22oi_1 _14302_ (.A1(_07976_),
    .A2(_08897_),
    .B1(_08898_),
    .B2(_07962_),
    .Y(_08899_));
 sky130_fd_sc_hd__mux2i_1 _14303_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .S(net3879),
    .Y(_08900_));
 sky130_fd_sc_hd__mux2i_1 _14304_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(net3879),
    .Y(_08901_));
 sky130_fd_sc_hd__a22oi_1 _14305_ (.A1(_07969_),
    .A2(_08900_),
    .B1(_08901_),
    .B2(_07983_),
    .Y(_08902_));
 sky130_fd_sc_hd__and3_4 _14306_ (.A(_07960_),
    .B(_08899_),
    .C(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__mux2_1 _14307_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net3867),
    .X(_08904_));
 sky130_fd_sc_hd__a221oi_1 _14308_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A2(_08829_),
    .B1(_08904_),
    .B2(net322),
    .C1(net3848),
    .Y(_08905_));
 sky130_fd_sc_hd__mux4_2 _14309_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S0(net3884),
    .S1(net3867),
    .X(_08906_));
 sky130_fd_sc_hd__nor2_1 _14310_ (.A(_07955_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nor4_1 _14311_ (.A(net3847),
    .B(net295),
    .C(_08905_),
    .D(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__mux4_2 _14312_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net3884),
    .S1(net3867),
    .X(_08909_));
 sky130_fd_sc_hd__nor2_4 _14313_ (.A(net3847),
    .B(net3849),
    .Y(_08910_));
 sky130_fd_sc_hd__mux4_2 _14314_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net3893),
    .S1(net3876),
    .X(_08911_));
 sky130_fd_sc_hd__a32oi_1 _14315_ (.A1(net294),
    .A2(_08909_),
    .A3(_08910_),
    .B1(net3798),
    .B2(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__mux4_2 _14316_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S0(net3893),
    .S1(net3876),
    .X(_08913_));
 sky130_fd_sc_hd__mux4_2 _14317_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S0(net3893),
    .S1(net3876),
    .X(_08914_));
 sky130_fd_sc_hd__a32oi_1 _14318_ (.A1(net294),
    .A2(_08820_),
    .A3(_08913_),
    .B1(_08914_),
    .B2(net351),
    .Y(_08915_));
 sky130_fd_sc_hd__nand2_1 _14319_ (.A(_08912_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__or3_4 _14320_ (.A(_08903_),
    .B(_08908_),
    .C(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1047 ();
 sky130_fd_sc_hd__a22o_4 _14322_ (.A1(net3840),
    .A2(_07912_),
    .B1(_08917_),
    .B2(_07888_),
    .X(_08919_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1046 ();
 sky130_fd_sc_hd__mux2_1 _14324_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .S(net3931),
    .X(_08921_));
 sky130_fd_sc_hd__nand2_1 _14325_ (.A(net3903),
    .B(_08921_),
    .Y(_08922_));
 sky130_fd_sc_hd__a211oi_1 _14326_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .A2(_08275_),
    .B1(net3899),
    .C1(net3913),
    .Y(_08923_));
 sky130_fd_sc_hd__mux2i_1 _14327_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S(net3931),
    .Y(_08924_));
 sky130_fd_sc_hd__mux2i_1 _14328_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net3931),
    .Y(_08925_));
 sky130_fd_sc_hd__a221oi_1 _14329_ (.A1(net413),
    .A2(_08924_),
    .B1(_08925_),
    .B2(_08282_),
    .C1(net3896),
    .Y(_08926_));
 sky130_fd_sc_hd__o2bb2ai_2 _14330_ (.A1_N(_08922_),
    .A2_N(_08923_),
    .B1(net3899),
    .B2(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__mux4_2 _14331_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S0(net3927),
    .S1(net3908),
    .X(_08928_));
 sky130_fd_sc_hd__mux4_2 _14332_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S0(net3927),
    .S1(net3908),
    .X(_08929_));
 sky130_fd_sc_hd__a22oi_2 _14333_ (.A1(_08126_),
    .A2(_08928_),
    .B1(_08929_),
    .B2(_08135_),
    .Y(_08930_));
 sky130_fd_sc_hd__mux4_2 _14334_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S0(net3931),
    .S1(net3913),
    .X(_08931_));
 sky130_fd_sc_hd__mux4_2 _14335_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net396),
    .S1(net3908),
    .X(_08932_));
 sky130_fd_sc_hd__mux4_2 _14336_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S0(net346),
    .S1(net3913),
    .X(_08933_));
 sky130_fd_sc_hd__a22o_1 _14337_ (.A1(_08126_),
    .A2(_08932_),
    .B1(_08933_),
    .B2(_08135_),
    .X(_08934_));
 sky130_fd_sc_hd__mux2i_1 _14338_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .S(net439),
    .Y(_08935_));
 sky130_fd_sc_hd__mux2i_1 _14339_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S(net439),
    .Y(_08936_));
 sky130_fd_sc_hd__o221ai_2 _14340_ (.A1(_08113_),
    .A2(_08935_),
    .B1(_08936_),
    .B2(_08119_),
    .C1(net3899),
    .Y(_08937_));
 sky130_fd_sc_hd__a211oi_2 _14341_ (.A1(_08111_),
    .A2(_08931_),
    .B1(_08934_),
    .C1(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__a21oi_4 _14342_ (.A1(_08927_),
    .A2(_08930_),
    .B1(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__nor2_1 _14343_ (.A(_08168_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__o22ai_1 _14344_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .B2(_08171_),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _14345_ (.A(_08172_),
    .B(_08917_),
    .Y(_08942_));
 sky130_fd_sc_hd__nor3_1 _14346_ (.A(_08940_),
    .B(_08941_),
    .C(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__o21ai_0 _14347_ (.A1(net3626),
    .A2(_08919_),
    .B1(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__xor2_1 _14348_ (.A(_08896_),
    .B(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__mux2i_2 _14349_ (.A0(_08939_),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .S(net293),
    .Y(_08946_));
 sky130_fd_sc_hd__o2bb2ai_4 _14350_ (.A1_N(\cs_registers_i.pc_id_i[8] ),
    .A2_N(_08202_),
    .B1(_08946_),
    .B2(net269),
    .Y(_08947_));
 sky130_fd_sc_hd__xnor2_1 _14351_ (.A(_08205_),
    .B(_08919_),
    .Y(_08948_));
 sky130_fd_sc_hd__xnor2_1 _14352_ (.A(net3615),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nor2_2 _14353_ (.A(net3755),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__a21oi_4 _14354_ (.A1(net3739),
    .A2(_08945_),
    .B1(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__nand2_2 _14355_ (.A(_08813_),
    .B(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__nand2_1 _14356_ (.A(_07857_),
    .B(_08896_),
    .Y(_08953_));
 sky130_fd_sc_hd__o21ai_1 _14357_ (.A1(_08316_),
    .A2(_08947_),
    .B1(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__or2_4 _14358_ (.A(_08804_),
    .B(_08812_),
    .X(_08955_));
 sky130_fd_sc_hd__nand2b_1 _14359_ (.A_N(_08943_),
    .B(_07857_),
    .Y(_08956_));
 sky130_fd_sc_hd__mux2i_1 _14360_ (.A0(_08205_),
    .A1(net291),
    .S(_08919_),
    .Y(_08957_));
 sky130_fd_sc_hd__a22o_1 _14361_ (.A1(net3593),
    .A2(_08955_),
    .B1(_08956_),
    .B2(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__o221ai_4 _14362_ (.A1(_08754_),
    .A2(_08952_),
    .B1(net3593),
    .B2(_08955_),
    .C1(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__xor2_1 _14363_ (.A(_08895_),
    .B(net327),
    .X(net180));
 sky130_fd_sc_hd__and2_4 _14364_ (.A(_08804_),
    .B(_08812_),
    .X(_08960_));
 sky130_fd_sc_hd__o21ai_2 _14365_ (.A1(net3541),
    .A2(_08960_),
    .B1(_08955_),
    .Y(_08961_));
 sky130_fd_sc_hd__xor2_1 _14366_ (.A(_08951_),
    .B(_08961_),
    .X(net179));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1044 ();
 sky130_fd_sc_hd__mux2_1 _14369_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .S(net3932),
    .X(_08964_));
 sky130_fd_sc_hd__a22oi_1 _14370_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .A2(_08275_),
    .B1(_08964_),
    .B2(net3904),
    .Y(_08965_));
 sky130_fd_sc_hd__mux4_2 _14371_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net3932),
    .S1(net3904),
    .X(_08966_));
 sky130_fd_sc_hd__nand2_1 _14372_ (.A(net3911),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__o211ai_1 _14373_ (.A1(net3911),
    .A2(_08965_),
    .B1(_08967_),
    .C1(net3781),
    .Y(_08968_));
 sky130_fd_sc_hd__mux4_2 _14374_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S0(net3930),
    .S1(net3911),
    .X(_08969_));
 sky130_fd_sc_hd__mux4_2 _14375_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S0(net3930),
    .S1(net3911),
    .X(_08970_));
 sky130_fd_sc_hd__o22a_1 _14376_ (.A1(net3770),
    .A2(_08969_),
    .B1(_08970_),
    .B2(_08389_),
    .X(_08971_));
 sky130_fd_sc_hd__mux4_2 _14377_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S0(net3927),
    .S1(net3911),
    .X(_08972_));
 sky130_fd_sc_hd__nand2_1 _14378_ (.A(net3904),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__mux4_2 _14379_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S0(net3927),
    .S1(net3911),
    .X(_08974_));
 sky130_fd_sc_hd__nand2_1 _14380_ (.A(_08109_),
    .B(_08974_),
    .Y(_08975_));
 sky130_fd_sc_hd__nand3_1 _14381_ (.A(net3774),
    .B(_08973_),
    .C(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__mux2_1 _14382_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .S(net3927),
    .X(_08977_));
 sky130_fd_sc_hd__nand2b_1 _14383_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .B(net3927),
    .Y(_08978_));
 sky130_fd_sc_hd__o221ai_1 _14384_ (.A1(net3927),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .B1(_08977_),
    .B2(net3911),
    .C1(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__mux2_1 _14385_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .S(net3927),
    .X(_08980_));
 sky130_fd_sc_hd__mux2_1 _14386_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S(net3927),
    .X(_08981_));
 sky130_fd_sc_hd__o211ai_1 _14387_ (.A1(net3911),
    .A2(_08980_),
    .B1(_08981_),
    .C1(net3904),
    .Y(_08982_));
 sky130_fd_sc_hd__a221oi_1 _14388_ (.A1(net3794),
    .A2(_08980_),
    .B1(_08977_),
    .B2(net3777),
    .C1(_08287_),
    .Y(_08983_));
 sky130_fd_sc_hd__o211ai_1 _14389_ (.A1(net3904),
    .A2(_08979_),
    .B1(_08982_),
    .C1(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand4_1 _14390_ (.A(_08968_),
    .B(_08971_),
    .C(_08976_),
    .D(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__inv_1 _14391_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .Y(_08986_));
 sky130_fd_sc_hd__mux2i_1 _14392_ (.A0(net3702),
    .A1(_08986_),
    .S(net3721),
    .Y(_08987_));
 sky130_fd_sc_hd__a22o_4 _14393_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(net3665),
    .B1(_08987_),
    .B2(net482),
    .X(_08988_));
 sky130_fd_sc_hd__mux2_1 _14394_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net3868),
    .X(_08989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1043 ();
 sky130_fd_sc_hd__a221oi_1 _14396_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .A2(net3764),
    .B1(_08989_),
    .B2(net322),
    .C1(net294),
    .Y(_08991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1042 ();
 sky130_fd_sc_hd__mux4_2 _14398_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net3884),
    .S1(net3868),
    .X(_08993_));
 sky130_fd_sc_hd__o21ai_0 _14399_ (.A1(_07927_),
    .A2(_08993_),
    .B1(_08910_),
    .Y(_08994_));
 sky130_fd_sc_hd__nor2_2 _14400_ (.A(_08991_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1040 ();
 sky130_fd_sc_hd__mux2i_1 _14403_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .S(net3871),
    .Y(_08998_));
 sky130_fd_sc_hd__mux2i_1 _14404_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S(net3871),
    .Y(_08999_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1039 ();
 sky130_fd_sc_hd__a22oi_1 _14406_ (.A1(net3806),
    .A2(_08998_),
    .B1(_08999_),
    .B2(net3811),
    .Y(_09001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1037 ();
 sky130_fd_sc_hd__mux2i_1 _14409_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(net3871),
    .Y(_09004_));
 sky130_fd_sc_hd__mux2i_1 _14410_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(net3871),
    .Y(_09005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1036 ();
 sky130_fd_sc_hd__a22oi_1 _14412_ (.A1(net3808),
    .A2(_09004_),
    .B1(_09005_),
    .B2(net3802),
    .Y(_09007_));
 sky130_fd_sc_hd__nand3_1 _14413_ (.A(net3765),
    .B(_09001_),
    .C(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__mux4_2 _14414_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09009_));
 sky130_fd_sc_hd__mux4_2 _14415_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09010_));
 sky130_fd_sc_hd__a22oi_2 _14416_ (.A1(net3801),
    .A2(_09009_),
    .B1(_09010_),
    .B2(net3798),
    .Y(_09011_));
 sky130_fd_sc_hd__mux2i_1 _14417_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S(net3871),
    .Y(_09012_));
 sky130_fd_sc_hd__mux2i_1 _14418_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .S(net3871),
    .Y(_09013_));
 sky130_fd_sc_hd__a22oi_1 _14419_ (.A1(net3811),
    .A2(_09012_),
    .B1(_09013_),
    .B2(net3808),
    .Y(_09014_));
 sky130_fd_sc_hd__mux2i_1 _14420_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .S(net3871),
    .Y(_09015_));
 sky130_fd_sc_hd__mux2i_1 _14421_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(net3871),
    .Y(_09016_));
 sky130_fd_sc_hd__a22oi_1 _14422_ (.A1(net3806),
    .A2(_09015_),
    .B1(_09016_),
    .B2(net3802),
    .Y(_09017_));
 sky130_fd_sc_hd__nand3_2 _14423_ (.A(net3752),
    .B(_09014_),
    .C(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand4b_1 _14424_ (.A_N(_08995_),
    .B(_09008_),
    .C(_09011_),
    .D(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__nor2_2 _14425_ (.A(_08348_),
    .B(net261),
    .Y(_09020_));
 sky130_fd_sc_hd__o31ai_1 _14426_ (.A1(_07892_),
    .A2(_07904_),
    .A3(_08352_),
    .B1(net3749),
    .Y(_09021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1035 ();
 sky130_fd_sc_hd__a22oi_1 _14428_ (.A1(net3836),
    .A2(_08355_),
    .B1(_09021_),
    .B2(net3895),
    .Y(_09023_));
 sky130_fd_sc_hd__nand3_1 _14429_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .B(_08632_),
    .C(_08355_),
    .Y(_09024_));
 sky130_fd_sc_hd__o221a_4 _14430_ (.A1(_08632_),
    .A2(_09023_),
    .B1(_09024_),
    .B2(net433),
    .C1(_08348_),
    .X(_09025_));
 sky130_fd_sc_hd__nor2_4 _14431_ (.A(_09020_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__xnor2_1 _14432_ (.A(net3626),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__xnor2_1 _14433_ (.A(_08988_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_2 _14434_ (.A(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B(_07864_),
    .Y(_09029_));
 sky130_fd_sc_hd__and4b_4 _14435_ (.A_N(_08995_),
    .B(_09008_),
    .C(_09011_),
    .D(_09018_),
    .X(_09030_));
 sky130_fd_sc_hd__o22ai_1 _14436_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .B2(_08171_),
    .Y(_09031_));
 sky130_fd_sc_hd__a221oi_2 _14437_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net3702),
    .B1(_09030_),
    .B2(net3736),
    .C1(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__o21ai_2 _14438_ (.A1(_09020_),
    .A2(_09025_),
    .B1(_08205_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_1 _14439_ (.A(_09032_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__xnor2_1 _14440_ (.A(_09029_),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__nor2_2 _14441_ (.A(net3747),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21oi_4 _14442_ (.A1(net3747),
    .A2(_09028_),
    .B1(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__nand2_8 _14443_ (.A(_07958_),
    .B(_07955_),
    .Y(_09038_));
 sky130_fd_sc_hd__mux4_2 _14444_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net3867),
    .S1(net3850),
    .X(_09039_));
 sky130_fd_sc_hd__mux2i_1 _14445_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .S(net3850),
    .Y(_09040_));
 sky130_fd_sc_hd__a21oi_1 _14446_ (.A1(net3850),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .B1(net3867),
    .Y(_09041_));
 sky130_fd_sc_hd__a211oi_1 _14447_ (.A1(net303),
    .A2(_09040_),
    .B1(_09041_),
    .C1(net322),
    .Y(_09042_));
 sky130_fd_sc_hd__a21oi_4 _14448_ (.A1(net3885),
    .A2(_09039_),
    .B1(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__mux2i_1 _14449_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .S(net3872),
    .Y(_09044_));
 sky130_fd_sc_hd__mux2i_1 _14450_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S(net3872),
    .Y(_09045_));
 sky130_fd_sc_hd__a22oi_1 _14451_ (.A1(net3804),
    .A2(_09044_),
    .B1(_09045_),
    .B2(net3809),
    .Y(_09046_));
 sky130_fd_sc_hd__mux2i_1 _14452_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S(net3872),
    .Y(_09047_));
 sky130_fd_sc_hd__mux2i_1 _14453_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(net3872),
    .Y(_09048_));
 sky130_fd_sc_hd__a22oi_1 _14454_ (.A1(net3811),
    .A2(_09047_),
    .B1(_09048_),
    .B2(net3803),
    .Y(_09049_));
 sky130_fd_sc_hd__mux4_2 _14455_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net3884),
    .S1(net3872),
    .X(_09050_));
 sky130_fd_sc_hd__mux4_2 _14456_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S0(net3884),
    .S1(net3872),
    .X(_09051_));
 sky130_fd_sc_hd__a22o_1 _14457_ (.A1(net3798),
    .A2(_09050_),
    .B1(_09051_),
    .B2(net276),
    .X(_09052_));
 sky130_fd_sc_hd__a31oi_1 _14458_ (.A1(net408),
    .A2(_09046_),
    .A3(_09049_),
    .B1(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__mux2i_1 _14459_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .S(net3872),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _14460_ (.A(net3809),
    .B(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__mux2i_1 _14461_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .S(net3872),
    .Y(_09056_));
 sky130_fd_sc_hd__mux2i_1 _14462_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S(net3872),
    .Y(_09057_));
 sky130_fd_sc_hd__a22oi_1 _14463_ (.A1(net3806),
    .A2(_09056_),
    .B1(_09057_),
    .B2(net3811),
    .Y(_09058_));
 sky130_fd_sc_hd__mux2i_1 _14464_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S(net3872),
    .Y(_09059_));
 sky130_fd_sc_hd__a21oi_1 _14465_ (.A1(net3803),
    .A2(_09059_),
    .B1(_08650_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand3_1 _14466_ (.A(_09055_),
    .B(_09058_),
    .C(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__o211ai_1 _14467_ (.A1(_09038_),
    .A2(_09043_),
    .B1(_09061_),
    .C1(_09053_),
    .Y(_09062_));
 sky130_fd_sc_hd__a22oi_1 _14468_ (.A1(net3837),
    .A2(_07912_),
    .B1(net3701),
    .B2(net3728),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_1 _14469_ (.A(_08205_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1033 ();
 sky130_fd_sc_hd__mux2i_1 _14472_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .S(net3930),
    .Y(_09067_));
 sky130_fd_sc_hd__mux2i_1 _14473_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .S(net3930),
    .Y(_09068_));
 sky130_fd_sc_hd__a22oi_1 _14474_ (.A1(net3777),
    .A2(_09067_),
    .B1(_09068_),
    .B2(net3794),
    .Y(_09069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1032 ();
 sky130_fd_sc_hd__mux2i_1 _14476_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S(net3930),
    .Y(_09071_));
 sky130_fd_sc_hd__mux2i_1 _14477_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S(net3930),
    .Y(_09072_));
 sky130_fd_sc_hd__a22oi_1 _14478_ (.A1(net3779),
    .A2(_09071_),
    .B1(_09072_),
    .B2(net3792),
    .Y(_09073_));
 sky130_fd_sc_hd__nand3_1 _14479_ (.A(_08694_),
    .B(_09069_),
    .C(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__mux4_2 _14480_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09075_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net3933),
    .X(_09076_));
 sky130_fd_sc_hd__a221o_1 _14482_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .A2(net3788),
    .B1(_09076_),
    .B2(net3914),
    .C1(net3901),
    .X(_09077_));
 sky130_fd_sc_hd__o211ai_1 _14483_ (.A1(_08109_),
    .A2(_09075_),
    .B1(_09077_),
    .C1(net3781),
    .Y(_09078_));
 sky130_fd_sc_hd__mux2i_1 _14484_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .S(net3930),
    .Y(_09079_));
 sky130_fd_sc_hd__mux2i_1 _14485_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .S(net3930),
    .Y(_09080_));
 sky130_fd_sc_hd__a22oi_1 _14486_ (.A1(net3777),
    .A2(_09079_),
    .B1(_09080_),
    .B2(net3794),
    .Y(_09081_));
 sky130_fd_sc_hd__mux2i_1 _14487_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S(net3930),
    .Y(_09082_));
 sky130_fd_sc_hd__mux2i_1 _14488_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S(net3930),
    .Y(_09083_));
 sky130_fd_sc_hd__a22oi_1 _14489_ (.A1(net3792),
    .A2(_09082_),
    .B1(_09083_),
    .B2(net3779),
    .Y(_09084_));
 sky130_fd_sc_hd__nand3_1 _14490_ (.A(net3773),
    .B(_09081_),
    .C(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__mux2i_1 _14491_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .S(net3930),
    .Y(_09086_));
 sky130_fd_sc_hd__mux2i_1 _14492_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S(net3930),
    .Y(_09087_));
 sky130_fd_sc_hd__a22oi_1 _14493_ (.A1(net3794),
    .A2(_09086_),
    .B1(_09087_),
    .B2(net3779),
    .Y(_09088_));
 sky130_fd_sc_hd__mux2i_1 _14494_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .S(net3930),
    .Y(_09089_));
 sky130_fd_sc_hd__mux2i_1 _14495_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(net3930),
    .Y(_09090_));
 sky130_fd_sc_hd__a22oi_1 _14496_ (.A1(net3777),
    .A2(_09089_),
    .B1(_09090_),
    .B2(net3792),
    .Y(_09091_));
 sky130_fd_sc_hd__nand3_1 _14497_ (.A(net3784),
    .B(_09088_),
    .C(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__and4_4 _14498_ (.A(_09078_),
    .B(_09074_),
    .C(_09085_),
    .D(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1030 ();
 sky130_fd_sc_hd__o22ai_1 _14501_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .B2(net3787),
    .Y(_09096_));
 sky130_fd_sc_hd__a21oi_1 _14502_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net400),
    .B1(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__o21ai_0 _14503_ (.A1(_08172_),
    .A2(net3701),
    .B1(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__nand2_1 _14504_ (.A(_07857_),
    .B(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__o211ai_1 _14505_ (.A1(_08442_),
    .A2(_09063_),
    .B1(_09064_),
    .C1(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1028 ();
 sky130_fd_sc_hd__nor2_1 _14508_ (.A(net3721),
    .B(net400),
    .Y(_09103_));
 sky130_fd_sc_hd__a21oi_1 _14509_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net3721),
    .B1(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1027 ();
 sky130_fd_sc_hd__nand2_1 _14511_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(net3665),
    .Y(_09106_));
 sky130_fd_sc_hd__o21ai_4 _14512_ (.A1(net3666),
    .A2(_09104_),
    .B1(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(net3744),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1026 ();
 sky130_fd_sc_hd__nand3_1 _14515_ (.A(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B(_08316_),
    .C(_07864_),
    .Y(_09110_));
 sky130_fd_sc_hd__nand2_2 _14516_ (.A(_09108_),
    .B(_09110_),
    .Y(_09111_));
 sky130_fd_sc_hd__xor2_1 _14517_ (.A(net3582),
    .B(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__and2_4 _14518_ (.A(_08895_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__o22ai_1 _14519_ (.A1(net300),
    .A2(_08845_),
    .B1(net474),
    .B2(net3744),
    .Y(_09114_));
 sky130_fd_sc_hd__a21o_1 _14520_ (.A1(net291),
    .A2(_08845_),
    .B1(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nor2_1 _14521_ (.A(_07857_),
    .B(_08890_),
    .Y(_09116_));
 sky130_fd_sc_hd__a21oi_1 _14522_ (.A1(_07857_),
    .A2(_08818_),
    .B1(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__a21oi_1 _14523_ (.A1(_09115_),
    .A2(_09117_),
    .B1(net3582),
    .Y(_09118_));
 sky130_fd_sc_hd__a31oi_1 _14524_ (.A1(net3582),
    .A2(_09115_),
    .A3(_09117_),
    .B1(_09111_),
    .Y(_09119_));
 sky130_fd_sc_hd__nor2_4 _14525_ (.A(_09118_),
    .B(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__a21oi_2 _14526_ (.A1(_08959_),
    .A2(_09113_),
    .B1(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__xnor2_4 _14527_ (.A(_09037_),
    .B(_09121_),
    .Y(net152));
 sky130_fd_sc_hd__a21oi_1 _14528_ (.A1(_08956_),
    .A2(_08957_),
    .B1(_08954_),
    .Y(_09122_));
 sky130_fd_sc_hd__maj3_2 _14529_ (.A(_09115_),
    .B(_09117_),
    .C(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__a31o_4 _14530_ (.A1(_08895_),
    .A2(_08951_),
    .A3(_08961_),
    .B1(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__xor2_4 _14531_ (.A(net3568),
    .B(_09124_),
    .X(net151));
 sky130_fd_sc_hd__mux2_1 _14532_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net3865),
    .X(_09125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1025 ();
 sky130_fd_sc_hd__a221oi_1 _14534_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .A2(net3764),
    .B1(_09125_),
    .B2(net3889),
    .C1(net3855),
    .Y(_09127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1024 ();
 sky130_fd_sc_hd__mux4_2 _14536_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net3889),
    .S1(net3865),
    .X(_09129_));
 sky130_fd_sc_hd__nor2_1 _14537_ (.A(_07927_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__mux2i_1 _14538_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(net3863),
    .Y(_09131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1023 ();
 sky130_fd_sc_hd__mux2i_1 _14540_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .S(net3863),
    .Y(_09133_));
 sky130_fd_sc_hd__a22oi_1 _14541_ (.A1(net3811),
    .A2(_09131_),
    .B1(_09133_),
    .B2(net3808),
    .Y(_09134_));
 sky130_fd_sc_hd__mux2i_1 _14542_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .S(net3863),
    .Y(_09135_));
 sky130_fd_sc_hd__mux2i_1 _14543_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S(net3863),
    .Y(_09136_));
 sky130_fd_sc_hd__a22oi_1 _14544_ (.A1(net3805),
    .A2(_09135_),
    .B1(_09136_),
    .B2(net3802),
    .Y(_09137_));
 sky130_fd_sc_hd__mux4_2 _14545_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net3883),
    .S1(net3863),
    .X(_09138_));
 sky130_fd_sc_hd__mux4_2 _14546_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net3883),
    .S1(net3863),
    .X(_09139_));
 sky130_fd_sc_hd__a22o_4 _14547_ (.A1(net3800),
    .A2(_09138_),
    .B1(_09139_),
    .B2(net3799),
    .X(_09140_));
 sky130_fd_sc_hd__a31oi_2 _14548_ (.A1(net3752),
    .A2(_09134_),
    .A3(_09137_),
    .B1(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__mux2i_1 _14549_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .S(net3863),
    .Y(_09142_));
 sky130_fd_sc_hd__mux2i_1 _14550_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S(net3863),
    .Y(_09143_));
 sky130_fd_sc_hd__a22oi_1 _14551_ (.A1(net3805),
    .A2(_09142_),
    .B1(_09143_),
    .B2(net3811),
    .Y(_09144_));
 sky130_fd_sc_hd__mux2i_1 _14552_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .S(net3863),
    .Y(_09145_));
 sky130_fd_sc_hd__mux2i_1 _14553_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(net3863),
    .Y(_09146_));
 sky130_fd_sc_hd__a22oi_2 _14554_ (.A1(net3808),
    .A2(_09145_),
    .B1(_09146_),
    .B2(net3802),
    .Y(_09147_));
 sky130_fd_sc_hd__nand3_1 _14555_ (.A(net3766),
    .B(_09144_),
    .C(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__o311a_4 _14556_ (.A1(_09038_),
    .A2(_09127_),
    .A3(_09130_),
    .B1(_09148_),
    .C1(_09141_),
    .X(_09149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1022 ();
 sky130_fd_sc_hd__a211oi_4 _14558_ (.A1(_07910_),
    .A2(_07908_),
    .B1(net3754),
    .C1(net3740),
    .Y(_09151_));
 sky130_fd_sc_hd__a21o_4 _14559_ (.A1(_07883_),
    .A2(_07886_),
    .B1(net3754),
    .X(_09152_));
 sky130_fd_sc_hd__a2111oi_4 _14560_ (.A1(_08352_),
    .A2(net3749),
    .B1(_08355_),
    .C1(_09152_),
    .D1(_07892_),
    .Y(_09153_));
 sky130_fd_sc_hd__or2_4 _14561_ (.A(_09151_),
    .B(net317),
    .X(_09154_));
 sky130_fd_sc_hd__nor2_2 _14562_ (.A(_07892_),
    .B(_08352_),
    .Y(_09155_));
 sky130_fd_sc_hd__o211a_4 _14563_ (.A1(net3740),
    .A2(_09155_),
    .B1(_08355_),
    .C1(net3836),
    .X(_09156_));
 sky130_fd_sc_hd__a211oi_2 _14564_ (.A1(net3939),
    .A2(_09154_),
    .B1(_09156_),
    .C1(_07888_),
    .Y(_09157_));
 sky130_fd_sc_hd__a21oi_4 _14565_ (.A1(_07888_),
    .A2(_09149_),
    .B1(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__mux2i_1 _14566_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .S(net3924),
    .Y(_09159_));
 sky130_fd_sc_hd__mux2i_1 _14567_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(net3924),
    .Y(_09160_));
 sky130_fd_sc_hd__a22oi_1 _14568_ (.A1(net3776),
    .A2(_09159_),
    .B1(_09160_),
    .B2(net3790),
    .Y(_09161_));
 sky130_fd_sc_hd__mux2i_1 _14569_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .S(net3924),
    .Y(_09162_));
 sky130_fd_sc_hd__mux2i_1 _14570_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S(net3924),
    .Y(_09163_));
 sky130_fd_sc_hd__a22oi_1 _14571_ (.A1(net3795),
    .A2(_09162_),
    .B1(_09163_),
    .B2(net3778),
    .Y(_09164_));
 sky130_fd_sc_hd__and3_4 _14572_ (.A(net3784),
    .B(_09161_),
    .C(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__mux2i_1 _14573_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(net3921),
    .Y(_09166_));
 sky130_fd_sc_hd__mux2i_1 _14574_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .S(net3921),
    .Y(_09167_));
 sky130_fd_sc_hd__a22oi_1 _14575_ (.A1(net3778),
    .A2(_09166_),
    .B1(_09167_),
    .B2(net3795),
    .Y(_09168_));
 sky130_fd_sc_hd__mux2i_1 _14576_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .S(net3921),
    .Y(_09169_));
 sky130_fd_sc_hd__mux2i_1 _14577_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S(net3921),
    .Y(_09170_));
 sky130_fd_sc_hd__a22oi_1 _14578_ (.A1(net3776),
    .A2(_09169_),
    .B1(_09170_),
    .B2(net3790),
    .Y(_09171_));
 sky130_fd_sc_hd__and3_4 _14579_ (.A(net3774),
    .B(_09168_),
    .C(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__mux2_1 _14580_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net3924),
    .X(_09173_));
 sky130_fd_sc_hd__a221oi_1 _14581_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .A2(net319),
    .B1(_09173_),
    .B2(net3910),
    .C1(net3905),
    .Y(_09174_));
 sky130_fd_sc_hd__mux4_2 _14582_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net3924),
    .S1(net3910),
    .X(_09175_));
 sky130_fd_sc_hd__o21ai_0 _14583_ (.A1(_08109_),
    .A2(_09175_),
    .B1(net3781),
    .Y(_09176_));
 sky130_fd_sc_hd__mux4_2 _14584_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09177_));
 sky130_fd_sc_hd__mux4_2 _14585_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09178_));
 sky130_fd_sc_hd__a22oi_2 _14586_ (.A1(_09177_),
    .A2(_08855_),
    .B1(_09178_),
    .B2(_08854_),
    .Y(_09179_));
 sky130_fd_sc_hd__o21ai_1 _14587_ (.A1(_09174_),
    .A2(_09176_),
    .B1(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__nor3_2 _14588_ (.A(_09165_),
    .B(_09172_),
    .C(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__o22ai_1 _14589_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .B2(net3786),
    .Y(_09182_));
 sky130_fd_sc_hd__a221oi_1 _14590_ (.A1(net3736),
    .A2(_09149_),
    .B1(net3699),
    .B2(net3949),
    .C1(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__o22ai_2 _14591_ (.A1(net3626),
    .A2(_09158_),
    .B1(_09183_),
    .B2(net3747),
    .Y(_09184_));
 sky130_fd_sc_hd__a21oi_4 _14592_ (.A1(net3624),
    .A2(_09158_),
    .B1(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__nor2_1 _14593_ (.A(net3723),
    .B(net3698),
    .Y(_09186_));
 sky130_fd_sc_hd__a21oi_1 _14594_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net3723),
    .B1(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__nand2_2 _14595_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(net3665),
    .Y(_09188_));
 sky130_fd_sc_hd__o21ai_4 _14596_ (.A1(net269),
    .A2(_09187_),
    .B1(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__and3_4 _14597_ (.A(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B(_07857_),
    .C(_07864_),
    .X(_09190_));
 sky130_fd_sc_hd__a21oi_4 _14598_ (.A1(net3745),
    .A2(_09189_),
    .B1(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__xor2_2 _14599_ (.A(_09185_),
    .B(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__nand2_8 _14600_ (.A(net3904),
    .B(_08694_),
    .Y(_09193_));
 sky130_fd_sc_hd__mux4_2 _14601_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net423),
    .S1(net3914),
    .X(_09194_));
 sky130_fd_sc_hd__mux4_2 _14602_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S0(net3929),
    .S1(net3914),
    .X(_09195_));
 sky130_fd_sc_hd__o22ai_1 _14603_ (.A1(_09193_),
    .A2(_09194_),
    .B1(_09195_),
    .B2(_08389_),
    .Y(_09196_));
 sky130_fd_sc_hd__mux4_2 _14604_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09197_));
 sky130_fd_sc_hd__nand2b_1 _14605_ (.A_N(_09197_),
    .B(net3901),
    .Y(_09198_));
 sky130_fd_sc_hd__mux2_1 _14606_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net3933),
    .X(_09199_));
 sky130_fd_sc_hd__a221o_1 _14607_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A2(net3788),
    .B1(_09199_),
    .B2(net3914),
    .C1(net3901),
    .X(_09200_));
 sky130_fd_sc_hd__a21oi_2 _14608_ (.A1(_09198_),
    .A2(_09200_),
    .B1(_08538_),
    .Y(_09201_));
 sky130_fd_sc_hd__mux4_2 _14609_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net3929),
    .S1(net3914),
    .X(_09202_));
 sky130_fd_sc_hd__mux4_2 _14610_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net424),
    .S1(net3914),
    .X(_09203_));
 sky130_fd_sc_hd__nand2_8 _14611_ (.A(_08109_),
    .B(net3772),
    .Y(_09204_));
 sky130_fd_sc_hd__o22ai_1 _14612_ (.A1(net3770),
    .A2(_09202_),
    .B1(_09203_),
    .B2(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand2_8 _14613_ (.A(_08109_),
    .B(_08694_),
    .Y(_09206_));
 sky130_fd_sc_hd__mux4_2 _14614_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net423),
    .S1(net3914),
    .X(_09207_));
 sky130_fd_sc_hd__mux4_2 _14615_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net424),
    .S1(net3914),
    .X(_09208_));
 sky130_fd_sc_hd__nand3b_1 _14616_ (.A_N(net3899),
    .B(net3903),
    .C(net3896),
    .Y(_09209_));
 sky130_fd_sc_hd__o22ai_1 _14617_ (.A1(_09206_),
    .A2(_09207_),
    .B1(_09208_),
    .B2(_09209_),
    .Y(_09210_));
 sky130_fd_sc_hd__or4_4 _14618_ (.A(_09196_),
    .B(_09205_),
    .C(_09201_),
    .D(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__inv_1 _14619_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .Y(_09212_));
 sky130_fd_sc_hd__mux2i_1 _14620_ (.A0(_09211_),
    .A1(_09212_),
    .S(net3721),
    .Y(_09213_));
 sky130_fd_sc_hd__a22o_4 _14621_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(net3665),
    .B1(_09213_),
    .B2(net482),
    .X(_09214_));
 sky130_fd_sc_hd__nand2_4 _14622_ (.A(net3745),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__nand3_2 _14623_ (.A(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .B(_07857_),
    .C(_07864_),
    .Y(_09216_));
 sky130_fd_sc_hd__nor2_1 _14624_ (.A(net3756),
    .B(_08988_),
    .Y(_09217_));
 sky130_fd_sc_hd__a21oi_2 _14625_ (.A1(net3756),
    .A2(_09029_),
    .B1(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__or2_4 _14626_ (.A(_09025_),
    .B(_09020_),
    .X(_09219_));
 sky130_fd_sc_hd__o221ai_4 _14627_ (.A1(net3747),
    .A2(_09032_),
    .B1(_09219_),
    .B2(_08442_),
    .C1(_09033_),
    .Y(_09220_));
 sky130_fd_sc_hd__maj3_1 _14628_ (.A(_09120_),
    .B(_09218_),
    .C(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__a31oi_4 _14629_ (.A1(net328),
    .A2(_09037_),
    .A3(_09113_),
    .B1(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand3_1 _14630_ (.A(_09215_),
    .B(_09216_),
    .C(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__o211ai_1 _14631_ (.A1(_09155_),
    .A2(net3740),
    .B1(_08355_),
    .C1(net3836),
    .Y(_09224_));
 sky130_fd_sc_hd__o21ai_2 _14632_ (.A1(_09151_),
    .A2(net317),
    .B1(net3944),
    .Y(_09225_));
 sky130_fd_sc_hd__mux4_2 _14633_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net3885),
    .S1(net3870),
    .X(_09226_));
 sky130_fd_sc_hd__mux4_2 _14634_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net3885),
    .S1(net3870),
    .X(_09227_));
 sky130_fd_sc_hd__mux2i_1 _14635_ (.A0(_09226_),
    .A1(_09227_),
    .S(net3817),
    .Y(_09228_));
 sky130_fd_sc_hd__mux2i_1 _14636_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .S(net3872),
    .Y(_09229_));
 sky130_fd_sc_hd__mux2i_1 _14637_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S(net3872),
    .Y(_09230_));
 sky130_fd_sc_hd__a22oi_1 _14638_ (.A1(net3809),
    .A2(_09229_),
    .B1(_09230_),
    .B2(net3811),
    .Y(_09231_));
 sky130_fd_sc_hd__mux2i_1 _14639_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .S(net3872),
    .Y(_09232_));
 sky130_fd_sc_hd__mux2i_1 _14640_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S(net3872),
    .Y(_09233_));
 sky130_fd_sc_hd__a22oi_1 _14641_ (.A1(net3804),
    .A2(_09232_),
    .B1(_09233_),
    .B2(net3803),
    .Y(_09234_));
 sky130_fd_sc_hd__mux4_2 _14642_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net3884),
    .S1(net3872),
    .X(_09235_));
 sky130_fd_sc_hd__mux4_2 _14643_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net3884),
    .S1(net3872),
    .X(_09236_));
 sky130_fd_sc_hd__a22o_1 _14644_ (.A1(net3801),
    .A2(_09235_),
    .B1(_09236_),
    .B2(net3798),
    .X(_09237_));
 sky130_fd_sc_hd__a31oi_2 _14645_ (.A1(net3765),
    .A2(_09231_),
    .A3(_09234_),
    .B1(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__mux4_2 _14646_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net3885),
    .S1(net303),
    .X(_09239_));
 sky130_fd_sc_hd__mux2_1 _14647_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net303),
    .X(_09240_));
 sky130_fd_sc_hd__a221o_1 _14648_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A2(net3764),
    .B1(_09240_),
    .B2(net3885),
    .C1(net295),
    .X(_09241_));
 sky130_fd_sc_hd__o211ai_1 _14649_ (.A1(net3817),
    .A2(_09239_),
    .B1(_09241_),
    .C1(net3762),
    .Y(_09242_));
 sky130_fd_sc_hd__o211a_4 _14650_ (.A1(_08650_),
    .A2(_09228_),
    .B1(_09238_),
    .C1(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__and2_4 _14651_ (.A(net3728),
    .B(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__a31oi_4 _14652_ (.A1(_08348_),
    .A2(net369),
    .A3(_09225_),
    .B1(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__o22ai_1 _14653_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .B2(_08171_),
    .Y(_09246_));
 sky130_fd_sc_hd__a221oi_1 _14654_ (.A1(net3949),
    .A2(_09211_),
    .B1(_09243_),
    .B2(net3736),
    .C1(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__o22ai_1 _14655_ (.A1(net3626),
    .A2(_09245_),
    .B1(_09247_),
    .B2(net3747),
    .Y(_09248_));
 sky130_fd_sc_hd__a21o_4 _14656_ (.A1(net3624),
    .A2(_09245_),
    .B1(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__a21oi_1 _14657_ (.A1(_09215_),
    .A2(_09216_),
    .B1(_09222_),
    .Y(_09250_));
 sky130_fd_sc_hd__a21oi_1 _14658_ (.A1(_09223_),
    .A2(_09249_),
    .B1(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__xor2_2 _14659_ (.A(_09192_),
    .B(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__inv_6 _14660_ (.A(net3498),
    .Y(net154));
 sky130_fd_sc_hd__nand2_4 _14661_ (.A(_09215_),
    .B(_09216_),
    .Y(_09253_));
 sky130_fd_sc_hd__xor2_2 _14662_ (.A(_09253_),
    .B(_09249_),
    .X(_09254_));
 sky130_fd_sc_hd__xnor2_4 _14663_ (.A(_09222_),
    .B(_09254_),
    .Y(net153));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1019 ();
 sky130_fd_sc_hd__mux4_2 _14667_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net3861),
    .S1(net3853),
    .X(_09258_));
 sky130_fd_sc_hd__mux4_2 _14668_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .S0(net3861),
    .S1(net3853),
    .X(_09259_));
 sky130_fd_sc_hd__mux2i_4 _14669_ (.A0(_09258_),
    .A1(_09259_),
    .S(_07935_),
    .Y(_09260_));
 sky130_fd_sc_hd__mux2i_1 _14670_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .S(net3866),
    .Y(_09261_));
 sky130_fd_sc_hd__mux2i_1 _14671_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S(net3866),
    .Y(_09262_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1018 ();
 sky130_fd_sc_hd__nand2_1 _14673_ (.A(net3866),
    .B(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .Y(_09264_));
 sky130_fd_sc_hd__mux2i_1 _14674_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net3866),
    .Y(_09265_));
 sky130_fd_sc_hd__mux4_2 _14675_ (.A0(_09261_),
    .A1(_09262_),
    .A2(_09264_),
    .A3(_09265_),
    .S0(net3891),
    .S1(_07927_),
    .X(_09266_));
 sky130_fd_sc_hd__mux2i_4 _14676_ (.A0(_09260_),
    .A1(_09266_),
    .S(_07958_),
    .Y(_09267_));
 sky130_fd_sc_hd__mux4_2 _14677_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net3861),
    .S1(net3853),
    .X(_09268_));
 sky130_fd_sc_hd__mux4_2 _14678_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .S0(net3861),
    .S1(net3853),
    .X(_09269_));
 sky130_fd_sc_hd__mux2_8 _14679_ (.A0(_09268_),
    .A1(_09269_),
    .S(_07935_),
    .X(_09270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1017 ();
 sky130_fd_sc_hd__mux4_2 _14681_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net3863),
    .S1(net3853),
    .X(_09272_));
 sky130_fd_sc_hd__mux4_2 _14682_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .S0(net3863),
    .S1(net3853),
    .X(_09273_));
 sky130_fd_sc_hd__mux2i_2 _14683_ (.A0(_09272_),
    .A1(_09273_),
    .S(_07935_),
    .Y(_09274_));
 sky130_fd_sc_hd__a2bb2oi_4 _14684_ (.A1_N(_08839_),
    .A2_N(_09270_),
    .B1(_09274_),
    .B2(net3766),
    .Y(_09275_));
 sky130_fd_sc_hd__o21ai_4 _14685_ (.A1(_09267_),
    .A2(net3849),
    .B1(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__a211oi_1 _14686_ (.A1(net3933),
    .A2(_09154_),
    .B1(_09156_),
    .C1(_07888_),
    .Y(_09277_));
 sky130_fd_sc_hd__a21oi_4 _14687_ (.A1(_07888_),
    .A2(net389),
    .B1(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1015 ();
 sky130_fd_sc_hd__mux4_2 _14690_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net3921),
    .S1(net3906),
    .X(_09281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1014 ();
 sky130_fd_sc_hd__mux4_2 _14692_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09283_));
 sky130_fd_sc_hd__o22ai_1 _14693_ (.A1(_08531_),
    .A2(_09281_),
    .B1(_09283_),
    .B2(net3769),
    .Y(_09284_));
 sky130_fd_sc_hd__nand2_1 _14694_ (.A(net283),
    .B(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1013 ();
 sky130_fd_sc_hd__mux4_2 _14696_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S0(net3921),
    .S1(net3906),
    .X(_09287_));
 sky130_fd_sc_hd__mux4_2 _14697_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09288_));
 sky130_fd_sc_hd__o22ai_1 _14698_ (.A1(_08531_),
    .A2(_09287_),
    .B1(_09288_),
    .B2(net3769),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _14699_ (.A(_08109_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1012 ();
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net3925),
    .X(_09292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1011 ();
 sky130_fd_sc_hd__a22oi_1 _14703_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .A2(net3789),
    .B1(_09292_),
    .B2(net3909),
    .Y(_09294_));
 sky130_fd_sc_hd__mux4_2 _14704_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net3925),
    .S1(net3909),
    .X(_09295_));
 sky130_fd_sc_hd__nand2_1 _14705_ (.A(net3902),
    .B(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__o211ai_1 _14706_ (.A1(net3902),
    .A2(_09294_),
    .B1(_09296_),
    .C1(net3781),
    .Y(_09297_));
 sky130_fd_sc_hd__mux4_2 _14707_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09298_));
 sky130_fd_sc_hd__mux4_2 _14708_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net3920),
    .S1(net3907),
    .X(_09299_));
 sky130_fd_sc_hd__mux2i_1 _14709_ (.A0(_09298_),
    .A1(_09299_),
    .S(_08109_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand2_1 _14710_ (.A(_08694_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand4_1 _14711_ (.A(_09285_),
    .B(_09290_),
    .C(_09297_),
    .D(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__o22ai_1 _14712_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .B2(net3786),
    .Y(_09303_));
 sky130_fd_sc_hd__a221oi_1 _14713_ (.A1(net3736),
    .A2(net389),
    .B1(net3697),
    .B2(net3949),
    .C1(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__o22ai_1 _14714_ (.A1(net3626),
    .A2(_09278_),
    .B1(_09304_),
    .B2(net3747),
    .Y(_09305_));
 sky130_fd_sc_hd__a21o_4 _14715_ (.A1(net3624),
    .A2(_09278_),
    .B1(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__nor2_1 _14716_ (.A(net3723),
    .B(net3697),
    .Y(_09307_));
 sky130_fd_sc_hd__a21oi_1 _14717_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net3723),
    .B1(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__nand2_1 _14718_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(net3665),
    .Y(_09309_));
 sky130_fd_sc_hd__o21ai_4 _14719_ (.A1(net269),
    .A2(_09308_),
    .B1(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__nand2_1 _14720_ (.A(net3737),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__nand3_1 _14721_ (.A(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B(net3739),
    .C(_07864_),
    .Y(_09312_));
 sky130_fd_sc_hd__nand2_2 _14722_ (.A(_09311_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__xor2_2 _14723_ (.A(_09306_),
    .B(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1010 ();
 sky130_fd_sc_hd__nand2_1 _14725_ (.A(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B(_07864_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_2 _14726_ (.A1(net315),
    .A2(net317),
    .B1(net3936),
    .Y(_09317_));
 sky130_fd_sc_hd__mux4_2 _14727_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net3889),
    .S1(net3875),
    .X(_09318_));
 sky130_fd_sc_hd__nor2_1 _14728_ (.A(_07927_),
    .B(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__mux2_1 _14729_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net3875),
    .X(_09320_));
 sky130_fd_sc_hd__a221oi_1 _14730_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .A2(net3764),
    .B1(_09320_),
    .B2(net3889),
    .C1(net3855),
    .Y(_09321_));
 sky130_fd_sc_hd__mux4_2 _14731_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net3883),
    .S1(net3865),
    .X(_09322_));
 sky130_fd_sc_hd__mux4_2 _14732_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net3883),
    .S1(net3865),
    .X(_09323_));
 sky130_fd_sc_hd__mux4_2 _14733_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net3883),
    .S1(net3863),
    .X(_09324_));
 sky130_fd_sc_hd__mux4_2 _14734_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net3883),
    .S1(net3863),
    .X(_09325_));
 sky130_fd_sc_hd__mux4_2 _14735_ (.A0(_09322_),
    .A1(_09323_),
    .A2(_09324_),
    .A3(_09325_),
    .S0(_07927_),
    .S1(net3844),
    .X(_09326_));
 sky130_fd_sc_hd__nand2_1 _14736_ (.A(net3848),
    .B(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__mux2i_1 _14737_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .S(net3863),
    .Y(_09328_));
 sky130_fd_sc_hd__mux2i_1 _14738_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(net3863),
    .Y(_09329_));
 sky130_fd_sc_hd__a22oi_1 _14739_ (.A1(net3805),
    .A2(_09328_),
    .B1(_09329_),
    .B2(net3811),
    .Y(_09330_));
 sky130_fd_sc_hd__mux2i_1 _14740_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .S(net3863),
    .Y(_09331_));
 sky130_fd_sc_hd__mux2i_1 _14741_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(net3863),
    .Y(_09332_));
 sky130_fd_sc_hd__a22oi_2 _14742_ (.A1(net3808),
    .A2(_09331_),
    .B1(_09332_),
    .B2(net3802),
    .Y(_09333_));
 sky130_fd_sc_hd__nand3_4 _14743_ (.A(net3752),
    .B(_09330_),
    .C(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__o311ai_2 _14744_ (.A1(_09038_),
    .A2(_09319_),
    .A3(_09321_),
    .B1(_09327_),
    .C1(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__nor2_2 _14745_ (.A(_08348_),
    .B(net3696),
    .Y(_09336_));
 sky130_fd_sc_hd__a31oi_4 _14746_ (.A1(_08348_),
    .A2(net369),
    .A3(_09317_),
    .B1(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__mux4_2 _14747_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net3921),
    .S1(net3906),
    .X(_09338_));
 sky130_fd_sc_hd__nand2_1 _14748_ (.A(net3905),
    .B(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__mux4_2 _14749_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net3921),
    .S1(net3906),
    .X(_09340_));
 sky130_fd_sc_hd__nand2_1 _14750_ (.A(_08109_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__a21oi_1 _14751_ (.A1(_09339_),
    .A2(_09341_),
    .B1(_08287_),
    .Y(_09342_));
 sky130_fd_sc_hd__mux4_2 _14752_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net3923),
    .S1(net3905),
    .X(_09343_));
 sky130_fd_sc_hd__nor2_1 _14753_ (.A(_08500_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__mux2_1 _14754_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .S(net3923),
    .X(_09345_));
 sky130_fd_sc_hd__a221oi_1 _14755_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .A2(_08275_),
    .B1(_09345_),
    .B2(net3905),
    .C1(net3910),
    .Y(_09346_));
 sky130_fd_sc_hd__nor3_2 _14756_ (.A(_08538_),
    .B(_09344_),
    .C(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__mux2i_1 _14757_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .S(net3921),
    .Y(_09348_));
 sky130_fd_sc_hd__mux2i_1 _14758_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(net3921),
    .Y(_09349_));
 sky130_fd_sc_hd__a22oi_1 _14759_ (.A1(net3776),
    .A2(_09348_),
    .B1(_09349_),
    .B2(net3790),
    .Y(_09350_));
 sky130_fd_sc_hd__mux2i_1 _14760_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .S(net3921),
    .Y(_09351_));
 sky130_fd_sc_hd__mux2i_1 _14761_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(net3921),
    .Y(_09352_));
 sky130_fd_sc_hd__a22oi_1 _14762_ (.A1(net3795),
    .A2(_09351_),
    .B1(_09352_),
    .B2(net3778),
    .Y(_09353_));
 sky130_fd_sc_hd__and3_4 _14763_ (.A(net3774),
    .B(_09350_),
    .C(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__mux2i_1 _14764_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S(net3923),
    .Y(_09355_));
 sky130_fd_sc_hd__mux2i_1 _14765_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .S(net3923),
    .Y(_09356_));
 sky130_fd_sc_hd__mux2i_1 _14766_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .S(net3923),
    .Y(_09357_));
 sky130_fd_sc_hd__a22o_1 _14767_ (.A1(net3776),
    .A2(_09356_),
    .B1(_09357_),
    .B2(net3795),
    .X(_09358_));
 sky130_fd_sc_hd__nor2b_1 _14768_ (.A(net3923),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .Y(_09359_));
 sky130_fd_sc_hd__a211oi_1 _14769_ (.A1(net3923),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .B1(_08266_),
    .C1(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__a2111oi_0 _14770_ (.A1(net3790),
    .A2(_09355_),
    .B1(_09358_),
    .C1(_09360_),
    .D1(_08531_),
    .Y(_09361_));
 sky130_fd_sc_hd__nor4_2 _14771_ (.A(_09342_),
    .B(_09347_),
    .C(_09354_),
    .D(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__o22ai_1 _14772_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .B2(_08171_),
    .Y(_09363_));
 sky130_fd_sc_hd__nor2_1 _14773_ (.A(_08172_),
    .B(net3696),
    .Y(_09364_));
 sky130_fd_sc_hd__a211oi_1 _14774_ (.A1(net3949),
    .A2(net3695),
    .B1(_09363_),
    .C1(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__o21ai_1 _14775_ (.A1(net3626),
    .A2(_09337_),
    .B1(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__xor2_1 _14776_ (.A(_09316_),
    .B(_09366_),
    .X(_09367_));
 sky130_fd_sc_hd__nor2_1 _14777_ (.A(net3721),
    .B(net3695),
    .Y(_09368_));
 sky130_fd_sc_hd__a21oi_1 _14778_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net3721),
    .B1(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__nand2_2 _14779_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(net3665),
    .Y(_09370_));
 sky130_fd_sc_hd__o21ai_4 _14780_ (.A1(net3666),
    .A2(_09369_),
    .B1(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _14781_ (.A(net3626),
    .B(_09337_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand2_2 _14782_ (.A(_09371_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__or2_0 _14783_ (.A(_09371_),
    .B(_09372_),
    .X(_09374_));
 sky130_fd_sc_hd__nand3_2 _14784_ (.A(net3747),
    .B(_09373_),
    .C(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__o21ai_4 _14785_ (.A1(net3737),
    .A2(_09367_),
    .B1(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand4_1 _14786_ (.A(_09037_),
    .B(_09192_),
    .C(_09254_),
    .D(_09376_),
    .Y(_09377_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1009 ();
 sky130_fd_sc_hd__nor2_1 _14788_ (.A(net3626),
    .B(_09337_),
    .Y(_09379_));
 sky130_fd_sc_hd__a211oi_1 _14789_ (.A1(net3626),
    .A2(_09337_),
    .B1(_09371_),
    .C1(net3756),
    .Y(_09380_));
 sky130_fd_sc_hd__a31oi_1 _14790_ (.A1(net3756),
    .A2(_09316_),
    .A3(_09365_),
    .B1(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand4_1 _14791_ (.A(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B(net3756),
    .C(_07864_),
    .D(_09366_),
    .Y(_09382_));
 sky130_fd_sc_hd__o21ai_2 _14792_ (.A1(net3756),
    .A2(_09373_),
    .B1(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand2_1 _14793_ (.A(_09185_),
    .B(_09191_),
    .Y(_09384_));
 sky130_fd_sc_hd__a31oi_1 _14794_ (.A1(_09253_),
    .A2(_09218_),
    .A3(_09220_),
    .B1(_09249_),
    .Y(_09385_));
 sky130_fd_sc_hd__a21oi_1 _14795_ (.A1(_09218_),
    .A2(_09220_),
    .B1(_09253_),
    .Y(_09386_));
 sky130_fd_sc_hd__o22ai_1 _14796_ (.A1(_09185_),
    .A2(_09191_),
    .B1(_09385_),
    .B2(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__and2_0 _14797_ (.A(_09384_),
    .B(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__o22ai_1 _14798_ (.A1(_09379_),
    .A2(_09381_),
    .B1(_09383_),
    .B2(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__o21ai_0 _14799_ (.A1(_09121_),
    .A2(_09377_),
    .B1(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__xor2_1 _14800_ (.A(_09314_),
    .B(_09390_),
    .X(net156));
 sky130_fd_sc_hd__inv_1 _14801_ (.A(_08960_),
    .Y(_09391_));
 sky130_fd_sc_hd__and4_4 _14802_ (.A(_09037_),
    .B(_09113_),
    .C(_09192_),
    .D(_09254_),
    .X(_09392_));
 sky130_fd_sc_hd__nand4b_1 _14803_ (.A_N(net3541),
    .B(_08951_),
    .C(_09391_),
    .D(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__maj3_1 _14804_ (.A(_09100_),
    .B(_09111_),
    .C(_09123_),
    .X(_09394_));
 sky130_fd_sc_hd__maj3_1 _14805_ (.A(_09218_),
    .B(_09220_),
    .C(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__maj3_1 _14806_ (.A(_09253_),
    .B(_09249_),
    .C(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__nor2_1 _14807_ (.A(_09185_),
    .B(_09191_),
    .Y(_09397_));
 sky130_fd_sc_hd__a21oi_2 _14808_ (.A1(_09384_),
    .A2(_09396_),
    .B1(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand3b_1 _14809_ (.A_N(_08955_),
    .B(_09392_),
    .C(_08951_),
    .Y(_09399_));
 sky130_fd_sc_hd__nand3_4 _14810_ (.A(_09393_),
    .B(_09398_),
    .C(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__xor2_2 _14811_ (.A(_09376_),
    .B(_09400_),
    .X(net155));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1008 ();
 sky130_fd_sc_hd__o21ai_2 _14813_ (.A1(net316),
    .A2(net317),
    .B1(net3901),
    .Y(_09402_));
 sky130_fd_sc_hd__mux4_2 _14814_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net322),
    .S1(net3866),
    .X(_09403_));
 sky130_fd_sc_hd__nand2_1 _14815_ (.A(net294),
    .B(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__mux4_2 _14816_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net322),
    .S1(net3866),
    .X(_09405_));
 sky130_fd_sc_hd__nand2_1 _14817_ (.A(net3817),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__and3_4 _14818_ (.A(net3848),
    .B(_09404_),
    .C(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__mux2_1 _14819_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .S(net294),
    .X(_09408_));
 sky130_fd_sc_hd__a22o_4 _14820_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .A2(net3815),
    .B1(_09408_),
    .B2(net262),
    .X(_09409_));
 sky130_fd_sc_hd__mux2i_1 _14821_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net303),
    .Y(_09410_));
 sky130_fd_sc_hd__mux2i_1 _14822_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S(net303),
    .Y(_09411_));
 sky130_fd_sc_hd__o221ai_2 _14823_ (.A1(net3814),
    .A2(_09410_),
    .B1(_09411_),
    .B2(_07951_),
    .C1(net3812),
    .Y(_09412_));
 sky130_fd_sc_hd__a21oi_4 _14824_ (.A1(_07935_),
    .A2(_09409_),
    .B1(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__mux2i_1 _14825_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S(net3864),
    .Y(_09414_));
 sky130_fd_sc_hd__mux2i_1 _14826_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .S(net3861),
    .Y(_09415_));
 sky130_fd_sc_hd__a22oi_2 _14827_ (.A1(net3810),
    .A2(_09414_),
    .B1(_09415_),
    .B2(net3809),
    .Y(_09416_));
 sky130_fd_sc_hd__mux2i_1 _14828_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .S(net3864),
    .Y(_09417_));
 sky130_fd_sc_hd__mux2i_1 _14829_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S(net3861),
    .Y(_09418_));
 sky130_fd_sc_hd__a22oi_1 _14830_ (.A1(net3804),
    .A2(_09417_),
    .B1(_09418_),
    .B2(net3803),
    .Y(_09419_));
 sky130_fd_sc_hd__mux4_2 _14831_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S0(net3882),
    .S1(net3861),
    .X(_09420_));
 sky130_fd_sc_hd__mux4_2 _14832_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S0(net3882),
    .S1(net3861),
    .X(_09421_));
 sky130_fd_sc_hd__a22o_4 _14833_ (.A1(net3799),
    .A2(_09420_),
    .B1(_09421_),
    .B2(net3800),
    .X(_09422_));
 sky130_fd_sc_hd__a31oi_4 _14834_ (.A1(net3751),
    .A2(_09416_),
    .A3(_09419_),
    .B1(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__o31ai_4 _14835_ (.A1(net3846),
    .A2(_09413_),
    .A3(_09407_),
    .B1(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_2 _14836_ (.A(net3718),
    .B(net410),
    .Y(_09425_));
 sky130_fd_sc_hd__a31oi_4 _14837_ (.A1(net3718),
    .A2(net3664),
    .A3(_09402_),
    .B1(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__mux2i_1 _14838_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .S(net346),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_1 _14839_ (.A(net260),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__mux2i_1 _14840_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S(net346),
    .Y(_09429_));
 sky130_fd_sc_hd__mux2i_1 _14841_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .S(net3919),
    .Y(_09430_));
 sky130_fd_sc_hd__a22oi_1 _14842_ (.A1(net3780),
    .A2(_09429_),
    .B1(_09430_),
    .B2(net3793),
    .Y(_09431_));
 sky130_fd_sc_hd__mux2i_1 _14843_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S(net3919),
    .Y(_09432_));
 sky130_fd_sc_hd__a21oi_1 _14844_ (.A1(_08147_),
    .A2(_09432_),
    .B1(net3769),
    .Y(_09433_));
 sky130_fd_sc_hd__nand3_4 _14845_ (.A(_09428_),
    .B(_09431_),
    .C(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__mux2i_1 _14846_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .S(net3919),
    .Y(_09435_));
 sky130_fd_sc_hd__mux2i_1 _14847_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .S(net3919),
    .Y(_09436_));
 sky130_fd_sc_hd__a22oi_1 _14848_ (.A1(net3793),
    .A2(_09435_),
    .B1(_09436_),
    .B2(net260),
    .Y(_09437_));
 sky130_fd_sc_hd__mux2i_1 _14849_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S(net3919),
    .Y(_09438_));
 sky130_fd_sc_hd__mux2i_1 _14850_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S(net3919),
    .Y(_09439_));
 sky130_fd_sc_hd__a22oi_1 _14851_ (.A1(net3780),
    .A2(_09438_),
    .B1(_09439_),
    .B2(net411),
    .Y(_09440_));
 sky130_fd_sc_hd__nand3_4 _14852_ (.A(_08694_),
    .B(_09437_),
    .C(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__mux4_2 _14853_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09442_));
 sky130_fd_sc_hd__nand2_1 _14854_ (.A(net3901),
    .B(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__a31oi_1 _14855_ (.A1(_08109_),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A3(net3788),
    .B1(net3897),
    .Y(_09444_));
 sky130_fd_sc_hd__mux2_1 _14856_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net439),
    .X(_09445_));
 sky130_fd_sc_hd__nand2_1 _14857_ (.A(net371),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__a31o_4 _14858_ (.A1(_09443_),
    .A2(_09444_),
    .A3(_09446_),
    .B1(net3896),
    .X(_09447_));
 sky130_fd_sc_hd__mux4_2 _14859_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .S0(net309),
    .S1(net3901),
    .X(_09448_));
 sky130_fd_sc_hd__nand2_1 _14860_ (.A(_08500_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__mux4_2 _14861_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net309),
    .S1(net3901),
    .X(_09450_));
 sky130_fd_sc_hd__a21oi_1 _14862_ (.A1(net3914),
    .A2(_09450_),
    .B1(net3768),
    .Y(_09451_));
 sky130_fd_sc_hd__a32oi_4 _14863_ (.A1(_09447_),
    .A2(_09441_),
    .A3(_09434_),
    .B1(_09449_),
    .B2(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__mux2i_1 _14864_ (.A0(net331),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .S(net3721),
    .Y(_09453_));
 sky130_fd_sc_hd__o2bb2ai_4 _14865_ (.A1_N(\cs_registers_i.pc_id_i[17] ),
    .A2_N(net3665),
    .B1(_09453_),
    .B2(net3666),
    .Y(_09454_));
 sky130_fd_sc_hd__xnor2_1 _14866_ (.A(net3626),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__xnor2_1 _14867_ (.A(_09426_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B(_07864_),
    .Y(_09457_));
 sky130_fd_sc_hd__nor2_1 _14869_ (.A(_08172_),
    .B(net409),
    .Y(_09458_));
 sky130_fd_sc_hd__o22ai_1 _14870_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .B2(_08171_),
    .Y(_09459_));
 sky130_fd_sc_hd__nor2_1 _14871_ (.A(_08168_),
    .B(net331),
    .Y(_09460_));
 sky130_fd_sc_hd__nor3_2 _14872_ (.A(_09458_),
    .B(_09459_),
    .C(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__o21ai_0 _14873_ (.A1(net3626),
    .A2(_09426_),
    .B1(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__xor2_1 _14874_ (.A(_09457_),
    .B(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__mux2i_4 _14875_ (.A0(_09456_),
    .A1(_09463_),
    .S(net3755),
    .Y(_09464_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1007 ();
 sky130_fd_sc_hd__nand2_1 _14877_ (.A(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B(_07864_),
    .Y(_09466_));
 sky130_fd_sc_hd__o21ai_2 _14878_ (.A1(net3700),
    .A2(net317),
    .B1(net3915),
    .Y(_09467_));
 sky130_fd_sc_hd__mux4_2 _14879_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net3885),
    .S1(net262),
    .X(_09468_));
 sky130_fd_sc_hd__nand2_1 _14880_ (.A(net294),
    .B(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__mux4_2 _14881_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net3885),
    .S1(net262),
    .X(_09470_));
 sky130_fd_sc_hd__nand2_2 _14882_ (.A(net3817),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand3_4 _14883_ (.A(net3848),
    .B(_09469_),
    .C(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__mux2_1 _14884_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .S(net295),
    .X(_09473_));
 sky130_fd_sc_hd__a22o_1 _14885_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .A2(net3816),
    .B1(_09473_),
    .B2(net262),
    .X(_09474_));
 sky130_fd_sc_hd__mux2i_1 _14886_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net262),
    .Y(_09475_));
 sky130_fd_sc_hd__mux2i_1 _14887_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(net262),
    .Y(_09476_));
 sky130_fd_sc_hd__o22ai_1 _14888_ (.A1(net3813),
    .A2(_09475_),
    .B1(_09476_),
    .B2(net430),
    .Y(_09477_));
 sky130_fd_sc_hd__a211o_4 _14889_ (.A1(_07935_),
    .A2(_09474_),
    .B1(_09477_),
    .C1(net3848),
    .X(_09478_));
 sky130_fd_sc_hd__mux2_1 _14890_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S(net3870),
    .X(_09479_));
 sky130_fd_sc_hd__mux2_1 _14891_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .S(net3871),
    .X(_09480_));
 sky130_fd_sc_hd__o22ai_2 _14892_ (.A1(net3813),
    .A2(_09479_),
    .B1(_09480_),
    .B2(_08570_),
    .Y(_09481_));
 sky130_fd_sc_hd__mux2i_1 _14893_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .S(net3870),
    .Y(_09482_));
 sky130_fd_sc_hd__mux2i_1 _14894_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(net3870),
    .Y(_09483_));
 sky130_fd_sc_hd__a22o_4 _14895_ (.A1(net3804),
    .A2(_09482_),
    .B1(_09483_),
    .B2(net3803),
    .X(_09484_));
 sky130_fd_sc_hd__mux4_2 _14896_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net322),
    .S1(net3872),
    .X(_09485_));
 sky130_fd_sc_hd__mux4_2 _14897_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net322),
    .S1(net3872),
    .X(_09486_));
 sky130_fd_sc_hd__a22oi_2 _14898_ (.A1(net3798),
    .A2(_09485_),
    .B1(_09486_),
    .B2(net3801),
    .Y(_09487_));
 sky130_fd_sc_hd__o31ai_4 _14899_ (.A1(_08650_),
    .A2(_09481_),
    .A3(_09484_),
    .B1(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__a31o_4 _14900_ (.A1(_07958_),
    .A2(_09472_),
    .A3(_09478_),
    .B1(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__nor2_2 _14901_ (.A(net3718),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__a31oi_4 _14902_ (.A1(net3718),
    .A2(net3664),
    .A3(_09467_),
    .B1(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .S(net3933),
    .X(_09492_));
 sky130_fd_sc_hd__a22oi_1 _14904_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .A2(_08275_),
    .B1(_09492_),
    .B2(net3901),
    .Y(_09493_));
 sky130_fd_sc_hd__mux4_2 _14905_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S0(net3933),
    .S1(net3901),
    .X(_09494_));
 sky130_fd_sc_hd__nand2_1 _14906_ (.A(net3914),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__o211ai_1 _14907_ (.A1(net3914),
    .A2(_09493_),
    .B1(_09495_),
    .C1(net3781),
    .Y(_09496_));
 sky130_fd_sc_hd__mux2_1 _14908_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .S(net309),
    .X(_09497_));
 sky130_fd_sc_hd__nand2b_1 _14909_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .B(net267),
    .Y(_09498_));
 sky130_fd_sc_hd__o221ai_1 _14910_ (.A1(net267),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .B1(_09497_),
    .B2(net3914),
    .C1(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__mux2_1 _14911_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .S(net309),
    .X(_09500_));
 sky130_fd_sc_hd__mux2_1 _14912_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(net309),
    .X(_09501_));
 sky130_fd_sc_hd__o211ai_1 _14913_ (.A1(net3914),
    .A2(_09500_),
    .B1(_09501_),
    .C1(net3901),
    .Y(_09502_));
 sky130_fd_sc_hd__a221oi_1 _14914_ (.A1(net3793),
    .A2(_09500_),
    .B1(_09497_),
    .B2(net3775),
    .C1(_08522_),
    .Y(_09503_));
 sky130_fd_sc_hd__o211ai_1 _14915_ (.A1(net3901),
    .A2(_09499_),
    .B1(_09502_),
    .C1(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__mux4_2 _14916_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net309),
    .S1(net3914),
    .X(_09505_));
 sky130_fd_sc_hd__mux4_2 _14917_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net309),
    .S1(net3914),
    .X(_09506_));
 sky130_fd_sc_hd__o22a_4 _14918_ (.A1(_09193_),
    .A2(_09505_),
    .B1(_09506_),
    .B2(_09206_),
    .X(_09507_));
 sky130_fd_sc_hd__mux4_2 _14919_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09508_));
 sky130_fd_sc_hd__mux4_2 _14920_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09509_));
 sky130_fd_sc_hd__o22a_1 _14921_ (.A1(net3770),
    .A2(_09508_),
    .B1(_09509_),
    .B2(_08389_),
    .X(_09510_));
 sky130_fd_sc_hd__nand4_1 _14922_ (.A(_09496_),
    .B(_09507_),
    .C(_09504_),
    .D(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__a31oi_4 _14923_ (.A1(_07958_),
    .A2(_09472_),
    .A3(_09478_),
    .B1(_09488_),
    .Y(_09512_));
 sky130_fd_sc_hd__o22ai_1 _14924_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .B2(_08171_),
    .Y(_09513_));
 sky130_fd_sc_hd__a221oi_2 _14925_ (.A1(net3949),
    .A2(net3693),
    .B1(_09512_),
    .B2(net3736),
    .C1(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21ai_0 _14926_ (.A1(net3626),
    .A2(_09491_),
    .B1(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__xor2_1 _14927_ (.A(_09466_),
    .B(_09515_),
    .X(_09516_));
 sky130_fd_sc_hd__nor2_1 _14928_ (.A(net3721),
    .B(net3693),
    .Y(_09517_));
 sky130_fd_sc_hd__a21oi_1 _14929_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net3722),
    .B1(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_2 _14930_ (.A(\cs_registers_i.pc_id_i[16] ),
    .B(net3665),
    .Y(_09519_));
 sky130_fd_sc_hd__o21ai_4 _14931_ (.A1(net3666),
    .A2(_09518_),
    .B1(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__xnor2_1 _14932_ (.A(_08205_),
    .B(_09491_),
    .Y(_09521_));
 sky130_fd_sc_hd__xnor2_1 _14933_ (.A(_09520_),
    .B(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand2_2 _14934_ (.A(net3745),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__o21ai_4 _14935_ (.A1(net3737),
    .A2(_09516_),
    .B1(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__nand2_1 _14936_ (.A(_09314_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__nor2_1 _14937_ (.A(_09377_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand3_1 _14938_ (.A(_09120_),
    .B(_09314_),
    .C(_09524_),
    .Y(_09527_));
 sky130_fd_sc_hd__nand2_1 _14939_ (.A(net3755),
    .B(_09466_),
    .Y(_09528_));
 sky130_fd_sc_hd__o21ai_2 _14940_ (.A1(net3739),
    .A2(_09520_),
    .B1(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__o22ai_1 _14941_ (.A1(net3745),
    .A2(_09514_),
    .B1(_09491_),
    .B2(net3626),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_2 _14942_ (.A1(net3624),
    .A2(_09491_),
    .B1(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand2_1 _14943_ (.A(_09529_),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__nor2_1 _14944_ (.A(_09529_),
    .B(_09531_),
    .Y(_09533_));
 sky130_fd_sc_hd__a31oi_1 _14945_ (.A1(_09306_),
    .A2(_09313_),
    .A3(_09532_),
    .B1(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__o221ai_1 _14946_ (.A1(_09389_),
    .A2(_09525_),
    .B1(_09527_),
    .B2(_09377_),
    .C1(_09534_),
    .Y(_09535_));
 sky130_fd_sc_hd__a31o_4 _14947_ (.A1(_09113_),
    .A2(_08959_),
    .A3(_09526_),
    .B1(_09535_),
    .X(_09536_));
 sky130_fd_sc_hd__xor2_4 _14948_ (.A(_09464_),
    .B(net419),
    .X(net158));
 sky130_fd_sc_hd__maj3_1 _14949_ (.A(_09306_),
    .B(_09313_),
    .C(_09383_),
    .X(_09537_));
 sky130_fd_sc_hd__a31oi_4 _14950_ (.A1(_09314_),
    .A2(_09376_),
    .A3(_09400_),
    .B1(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__xnor2_2 _14951_ (.A(_09524_),
    .B(_09538_),
    .Y(net157));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1006 ();
 sky130_fd_sc_hd__nand2_1 _14953_ (.A(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B(_07864_),
    .Y(_09540_));
 sky130_fd_sc_hd__a21oi_4 _14954_ (.A1(net3896),
    .A2(_09154_),
    .B1(_09156_),
    .Y(_09541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1005 ();
 sky130_fd_sc_hd__mux4_2 _14956_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net322),
    .S1(net3866),
    .X(_09543_));
 sky130_fd_sc_hd__nand2_1 _14957_ (.A(net294),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__mux4_2 _14958_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net3887),
    .S1(net3866),
    .X(_09545_));
 sky130_fd_sc_hd__nand2_1 _14959_ (.A(_07927_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__and3_4 _14960_ (.A(net3848),
    .B(_09544_),
    .C(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__mux2_1 _14961_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .S(net295),
    .X(_09548_));
 sky130_fd_sc_hd__a22o_1 _14962_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .A2(net3815),
    .B1(_09548_),
    .B2(net262),
    .X(_09549_));
 sky130_fd_sc_hd__mux2i_1 _14963_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net303),
    .Y(_09550_));
 sky130_fd_sc_hd__mux2i_1 _14964_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S(net303),
    .Y(_09551_));
 sky130_fd_sc_hd__o221ai_1 _14965_ (.A1(net3814),
    .A2(_09550_),
    .B1(_09551_),
    .B2(net430),
    .C1(net3812),
    .Y(_09552_));
 sky130_fd_sc_hd__a21oi_2 _14966_ (.A1(_07935_),
    .A2(_09549_),
    .B1(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__mux2i_1 _14967_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S(net3861),
    .Y(_09554_));
 sky130_fd_sc_hd__mux2i_1 _14968_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .S(net3861),
    .Y(_09555_));
 sky130_fd_sc_hd__a22oi_2 _14969_ (.A1(net3810),
    .A2(_09554_),
    .B1(_09555_),
    .B2(net3809),
    .Y(_09556_));
 sky130_fd_sc_hd__mux2i_1 _14970_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .S(net3861),
    .Y(_09557_));
 sky130_fd_sc_hd__mux2i_1 _14971_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S(net3861),
    .Y(_09558_));
 sky130_fd_sc_hd__a22oi_2 _14972_ (.A1(net3804),
    .A2(_09557_),
    .B1(_09558_),
    .B2(net3803),
    .Y(_09559_));
 sky130_fd_sc_hd__mux4_2 _14973_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net3881),
    .S1(net3861),
    .X(_09560_));
 sky130_fd_sc_hd__mux4_2 _14974_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net3881),
    .S1(net3861),
    .X(_09561_));
 sky130_fd_sc_hd__a22o_4 _14975_ (.A1(net3800),
    .A2(_09560_),
    .B1(_09561_),
    .B2(net3799),
    .X(_09562_));
 sky130_fd_sc_hd__a31oi_4 _14976_ (.A1(net3751),
    .A2(_09556_),
    .A3(_09559_),
    .B1(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__o31ai_4 _14977_ (.A1(net3844),
    .A2(_09553_),
    .A3(_09547_),
    .B1(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__nand2_1 _14978_ (.A(net3728),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__o21ai_4 _14979_ (.A1(net3728),
    .A2(_09541_),
    .B1(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__mux2i_1 _14980_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S(net3933),
    .Y(_09567_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_08261_),
    .B(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__mux2i_1 _14982_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net3933),
    .Y(_09569_));
 sky130_fd_sc_hd__mux2i_1 _14983_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .S(net3933),
    .Y(_09570_));
 sky130_fd_sc_hd__o22ai_1 _14984_ (.A1(_08266_),
    .A2(_09569_),
    .B1(_09570_),
    .B2(_08374_),
    .Y(_09571_));
 sky130_fd_sc_hd__a2111oi_4 _14985_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A2(net3767),
    .B1(_09568_),
    .C1(_09571_),
    .D1(_08538_),
    .Y(_09572_));
 sky130_fd_sc_hd__inv_6 _14986_ (.A(net3896),
    .Y(_09573_));
 sky130_fd_sc_hd__mux4_2 _14987_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09574_));
 sky130_fd_sc_hd__mux4_2 _14988_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09575_));
 sky130_fd_sc_hd__mux4_2 _14989_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09576_));
 sky130_fd_sc_hd__mux4_2 _14990_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09577_));
 sky130_fd_sc_hd__mux4_2 _14991_ (.A0(_09574_),
    .A1(_09575_),
    .A2(_09576_),
    .A3(_09577_),
    .S0(_08109_),
    .S1(net3898),
    .X(_09578_));
 sky130_fd_sc_hd__mux4_2 _14992_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net309),
    .S1(net3914),
    .X(_09579_));
 sky130_fd_sc_hd__mux4_2 _14993_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net267),
    .S1(net3913),
    .X(_09580_));
 sky130_fd_sc_hd__mux2_4 _14994_ (.A0(_09579_),
    .A1(_09580_),
    .S(_08109_),
    .X(_09581_));
 sky130_fd_sc_hd__o22ai_4 _14995_ (.A1(_09578_),
    .A2(_09573_),
    .B1(_09581_),
    .B2(net3768),
    .Y(_09582_));
 sky130_fd_sc_hd__nor2_4 _14996_ (.A(_09582_),
    .B(_09572_),
    .Y(_09583_));
 sky130_fd_sc_hd__nor2_1 _14997_ (.A(_08168_),
    .B(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__nor2_1 _14998_ (.A(_08172_),
    .B(_09564_),
    .Y(_09585_));
 sky130_fd_sc_hd__o22ai_1 _14999_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .B2(_08171_),
    .Y(_09586_));
 sky130_fd_sc_hd__nor3_2 _15000_ (.A(_09584_),
    .B(_09585_),
    .C(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__o21ai_0 _15001_ (.A1(net3626),
    .A2(_09566_),
    .B1(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__xor2_1 _15002_ (.A(_09540_),
    .B(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1004 ();
 sky130_fd_sc_hd__mux2i_2 _15004_ (.A0(_09583_),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .S(net3721),
    .Y(_09591_));
 sky130_fd_sc_hd__nand2_1 _15005_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(net3665),
    .Y(_09592_));
 sky130_fd_sc_hd__o21ai_4 _15006_ (.A1(net3666),
    .A2(_09591_),
    .B1(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__xnor2_1 _15007_ (.A(_08205_),
    .B(_09566_),
    .Y(_09594_));
 sky130_fd_sc_hd__xnor2_1 _15008_ (.A(_09593_),
    .B(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand2_2 _15009_ (.A(net3745),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__o21ai_4 _15010_ (.A1(net3745),
    .A2(_09589_),
    .B1(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__o21ai_4 _15011_ (.A1(net3700),
    .A2(net317),
    .B1(net3897),
    .Y(_09598_));
 sky130_fd_sc_hd__mux4_2 _15012_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09599_));
 sky130_fd_sc_hd__nand2_1 _15013_ (.A(net295),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__mux4_2 _15014_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09601_));
 sky130_fd_sc_hd__nand2_1 _15015_ (.A(_07927_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__and3_4 _15016_ (.A(net3849),
    .B(_09600_),
    .C(_09602_),
    .X(_09603_));
 sky130_fd_sc_hd__mux2_1 _15017_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .S(net3850),
    .X(_09604_));
 sky130_fd_sc_hd__a22o_1 _15018_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .A2(net3816),
    .B1(_09604_),
    .B2(net3871),
    .X(_09605_));
 sky130_fd_sc_hd__mux2i_1 _15019_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net3871),
    .Y(_09606_));
 sky130_fd_sc_hd__mux2i_1 _15020_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S(net3871),
    .Y(_09607_));
 sky130_fd_sc_hd__o221ai_1 _15021_ (.A1(net365),
    .A2(_09606_),
    .B1(_09607_),
    .B2(net427),
    .C1(_07955_),
    .Y(_09608_));
 sky130_fd_sc_hd__a21oi_2 _15022_ (.A1(_07935_),
    .A2(_09605_),
    .B1(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__mux2i_1 _15023_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S(net3871),
    .Y(_09610_));
 sky130_fd_sc_hd__mux2i_1 _15024_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .S(net3871),
    .Y(_09611_));
 sky130_fd_sc_hd__a22oi_2 _15025_ (.A1(net3811),
    .A2(_09610_),
    .B1(_09611_),
    .B2(net3808),
    .Y(_09612_));
 sky130_fd_sc_hd__mux2i_1 _15026_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .S(net3871),
    .Y(_09613_));
 sky130_fd_sc_hd__mux2i_1 _15027_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S(net3871),
    .Y(_09614_));
 sky130_fd_sc_hd__a22oi_2 _15028_ (.A1(net3806),
    .A2(_09613_),
    .B1(_09614_),
    .B2(net3802),
    .Y(_09615_));
 sky130_fd_sc_hd__mux4_2 _15029_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09616_));
 sky130_fd_sc_hd__mux4_2 _15030_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net3884),
    .S1(net3868),
    .X(_09617_));
 sky130_fd_sc_hd__a22o_4 _15031_ (.A1(net3798),
    .A2(_09616_),
    .B1(_09617_),
    .B2(net3801),
    .X(_09618_));
 sky130_fd_sc_hd__a31oi_4 _15032_ (.A1(net3752),
    .A2(_09612_),
    .A3(_09615_),
    .B1(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__o31ai_4 _15033_ (.A1(net3847),
    .A2(_09603_),
    .A3(_09609_),
    .B1(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__nor2_1 _15034_ (.A(_08348_),
    .B(net3692),
    .Y(_09621_));
 sky130_fd_sc_hd__a31oi_4 _15035_ (.A1(_08348_),
    .A2(net3664),
    .A3(_09598_),
    .B1(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nor2_2 _15036_ (.A(net3626),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__nor2_1 _15037_ (.A(_08172_),
    .B(net3692),
    .Y(_09624_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1002 ();
 sky130_fd_sc_hd__o22ai_1 _15040_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .B2(net3786),
    .Y(_09627_));
 sky130_fd_sc_hd__nor2_1 _15041_ (.A(_09624_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__mux2i_1 _15042_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S(net267),
    .Y(_09629_));
 sky130_fd_sc_hd__mux2i_1 _15043_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .S(net267),
    .Y(_09630_));
 sky130_fd_sc_hd__o22ai_1 _15044_ (.A1(net3783),
    .A2(_09629_),
    .B1(_09630_),
    .B2(net3771),
    .Y(_09631_));
 sky130_fd_sc_hd__mux2i_1 _15045_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net267),
    .Y(_09632_));
 sky130_fd_sc_hd__o2bb2ai_1 _15046_ (.A1_N(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .A2_N(net3767),
    .B1(_09632_),
    .B2(net3782),
    .Y(_09633_));
 sky130_fd_sc_hd__nor3_2 _15047_ (.A(_08538_),
    .B(_09631_),
    .C(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__mux2_1 _15048_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .S(net3927),
    .X(_09635_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .S(net3927),
    .X(_09636_));
 sky130_fd_sc_hd__a221oi_1 _15050_ (.A1(net3794),
    .A2(_09635_),
    .B1(_09636_),
    .B2(net3777),
    .C1(_08287_),
    .Y(_09637_));
 sky130_fd_sc_hd__mux2_1 _15051_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S(net3927),
    .X(_09638_));
 sky130_fd_sc_hd__o211ai_1 _15052_ (.A1(net3911),
    .A2(_09635_),
    .B1(_09638_),
    .C1(net3904),
    .Y(_09639_));
 sky130_fd_sc_hd__mux2_1 _15053_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S(net3927),
    .X(_09640_));
 sky130_fd_sc_hd__o211ai_1 _15054_ (.A1(net3911),
    .A2(_09636_),
    .B1(_09640_),
    .C1(_08109_),
    .Y(_09641_));
 sky130_fd_sc_hd__and3_4 _15055_ (.A(_09637_),
    .B(_09639_),
    .C(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__nor2_2 _15056_ (.A(_09634_),
    .B(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__mux4_2 _15057_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net3927),
    .S1(net3911),
    .X(_09644_));
 sky130_fd_sc_hd__mux4_2 _15058_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net3930),
    .S1(net3911),
    .X(_09645_));
 sky130_fd_sc_hd__o22ai_1 _15059_ (.A1(net3770),
    .A2(_09644_),
    .B1(_09645_),
    .B2(_08389_),
    .Y(_09646_));
 sky130_fd_sc_hd__mux4_2 _15060_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S0(net3927),
    .S1(net3911),
    .X(_09647_));
 sky130_fd_sc_hd__nor3_2 _15061_ (.A(net3904),
    .B(_08522_),
    .C(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__mux4_2 _15062_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S0(net3927),
    .S1(net3911),
    .X(_09649_));
 sky130_fd_sc_hd__nor2_1 _15063_ (.A(_09209_),
    .B(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__nor3_4 _15064_ (.A(_09646_),
    .B(_09648_),
    .C(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_8 _15065_ (.A(_09643_),
    .B(net3735),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_1 _15066_ (.A(net3949),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21oi_2 _15067_ (.A1(_09628_),
    .A2(_09653_),
    .B1(net3745),
    .Y(_09654_));
 sky130_fd_sc_hd__a211oi_4 _15068_ (.A1(net3624),
    .A2(_09622_),
    .B1(_09623_),
    .C1(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nor2_2 _15069_ (.A(net3626),
    .B(_09426_),
    .Y(_09656_));
 sky130_fd_sc_hd__nor2_1 _15070_ (.A(net3745),
    .B(_09461_),
    .Y(_09657_));
 sky130_fd_sc_hd__a211oi_4 _15071_ (.A1(net3624),
    .A2(_09426_),
    .B1(_09656_),
    .C1(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand2_1 _15072_ (.A(net3755),
    .B(_09457_),
    .Y(_09659_));
 sky130_fd_sc_hd__o21ai_4 _15073_ (.A1(net3739),
    .A2(_09454_),
    .B1(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__nand2_1 _15074_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .B(net3721),
    .Y(_09661_));
 sky130_fd_sc_hd__o21ai_0 _15075_ (.A1(net3721),
    .A2(_09652_),
    .B1(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__a22o_4 _15076_ (.A1(\cs_registers_i.pc_id_i[18] ),
    .A2(net3665),
    .B1(_09662_),
    .B2(net482),
    .X(_09663_));
 sky130_fd_sc_hd__and3_1 _15077_ (.A(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B(net3755),
    .C(_07864_),
    .X(_09664_));
 sky130_fd_sc_hd__a21oi_2 _15078_ (.A1(net3745),
    .A2(_09663_),
    .B1(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__o31ai_2 _15079_ (.A1(_09655_),
    .A2(_09658_),
    .A3(_09660_),
    .B1(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o21ai_2 _15080_ (.A1(_09658_),
    .A2(_09660_),
    .B1(_09655_),
    .Y(_09667_));
 sky130_fd_sc_hd__xor2_1 _15081_ (.A(_09665_),
    .B(_09655_),
    .X(_09668_));
 sky130_fd_sc_hd__and2_4 _15082_ (.A(_09464_),
    .B(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__a22o_4 _15083_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_09669_),
    .B2(_09536_),
    .X(_09670_));
 sky130_fd_sc_hd__xor2_4 _15084_ (.A(_09597_),
    .B(_09670_),
    .X(net160));
 sky130_fd_sc_hd__nand2_1 _15085_ (.A(_09464_),
    .B(_09524_),
    .Y(_09671_));
 sky130_fd_sc_hd__or2_0 _15086_ (.A(_09529_),
    .B(_09531_),
    .X(_09672_));
 sky130_fd_sc_hd__maj3_1 _15087_ (.A(_09672_),
    .B(_09658_),
    .C(_09660_),
    .X(_09673_));
 sky130_fd_sc_hd__o21ai_0 _15088_ (.A1(_09538_),
    .A2(_09671_),
    .B1(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__xnor2_1 _15089_ (.A(_09668_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__inv_1 _15090_ (.A(net3497),
    .Y(net159));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1001 ();
 sky130_fd_sc_hd__nand2_2 _15092_ (.A(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B(_07864_),
    .Y(_09677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_999 ();
 sky130_fd_sc_hd__nor3b_4 _15095_ (.A(_07911_),
    .B(net3754),
    .C_N(net3836),
    .Y(_09680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_998 ();
 sky130_fd_sc_hd__a21oi_4 _15097_ (.A1(net3858),
    .A2(net3700),
    .B1(_09680_),
    .Y(_09682_));
 sky130_fd_sc_hd__mux4_2 _15098_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net3893),
    .S1(net3878),
    .X(_09683_));
 sky130_fd_sc_hd__nand2_1 _15099_ (.A(net3854),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__mux4_2 _15100_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net3893),
    .S1(net3878),
    .X(_09685_));
 sky130_fd_sc_hd__nand2_1 _15101_ (.A(_07927_),
    .B(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__and3_4 _15102_ (.A(net3849),
    .B(_09684_),
    .C(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__mux2_1 _15103_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .S(net3850),
    .X(_09688_));
 sky130_fd_sc_hd__a22o_1 _15104_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .A2(net345),
    .B1(_09688_),
    .B2(net3868),
    .X(_09689_));
 sky130_fd_sc_hd__mux2i_1 _15105_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net303),
    .Y(_09690_));
 sky130_fd_sc_hd__mux2i_1 _15106_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S(net303),
    .Y(_09691_));
 sky130_fd_sc_hd__o221ai_1 _15107_ (.A1(_07945_),
    .A2(_09690_),
    .B1(_09691_),
    .B2(_07951_),
    .C1(_07955_),
    .Y(_09692_));
 sky130_fd_sc_hd__a21oi_1 _15108_ (.A1(_07935_),
    .A2(_09689_),
    .B1(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__mux2i_1 _15109_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S(net3878),
    .Y(_09694_));
 sky130_fd_sc_hd__mux2i_1 _15110_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .S(net3878),
    .Y(_09695_));
 sky130_fd_sc_hd__a22oi_1 _15111_ (.A1(net3811),
    .A2(_09694_),
    .B1(_09695_),
    .B2(net3808),
    .Y(_09696_));
 sky130_fd_sc_hd__mux2i_1 _15112_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .S(net3878),
    .Y(_09697_));
 sky130_fd_sc_hd__mux2i_1 _15113_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S(net3878),
    .Y(_09698_));
 sky130_fd_sc_hd__a22oi_1 _15114_ (.A1(net3806),
    .A2(_09697_),
    .B1(_09698_),
    .B2(net3802),
    .Y(_09699_));
 sky130_fd_sc_hd__mux4_2 _15115_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S0(net3893),
    .S1(net3878),
    .X(_09700_));
 sky130_fd_sc_hd__mux4_2 _15116_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net3893),
    .S1(net3878),
    .X(_09701_));
 sky130_fd_sc_hd__a22o_4 _15117_ (.A1(net351),
    .A2(_09700_),
    .B1(_09701_),
    .B2(net3798),
    .X(_09702_));
 sky130_fd_sc_hd__a31oi_4 _15118_ (.A1(net3752),
    .A2(_09696_),
    .A3(_09699_),
    .B1(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__o31ai_4 _15119_ (.A1(net3847),
    .A2(_09687_),
    .A3(_09693_),
    .B1(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(net3728),
    .B(net3691),
    .Y(_09705_));
 sky130_fd_sc_hd__o21ai_4 _15121_ (.A1(net3728),
    .A2(_09682_),
    .B1(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__mux4_2 _15122_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09707_));
 sky130_fd_sc_hd__mux4_2 _15123_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09708_));
 sky130_fd_sc_hd__mux4_2 _15124_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09709_));
 sky130_fd_sc_hd__mux4_2 _15125_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09710_));
 sky130_fd_sc_hd__mux4_2 _15126_ (.A0(_09707_),
    .A1(_09708_),
    .A2(_09709_),
    .A3(_09710_),
    .S0(net3903),
    .S1(net3899),
    .X(_09711_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .S(net3931),
    .X(_09712_));
 sky130_fd_sc_hd__mux2_1 _15128_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S(net3931),
    .X(_09713_));
 sky130_fd_sc_hd__mux2_1 _15129_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net3931),
    .X(_09714_));
 sky130_fd_sc_hd__a222oi_1 _15130_ (.A1(net263),
    .A2(_09712_),
    .B1(_09713_),
    .B2(net3792),
    .C1(_09714_),
    .C2(net3779),
    .Y(_09715_));
 sky130_fd_sc_hd__a21oi_2 _15131_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A2(net3767),
    .B1(_08538_),
    .Y(_09716_));
 sky130_fd_sc_hd__mux4_2 _15132_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09717_));
 sky130_fd_sc_hd__mux4_2 _15133_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net3926),
    .S1(net3912),
    .X(_09718_));
 sky130_fd_sc_hd__o22ai_2 _15134_ (.A1(net3770),
    .A2(_09717_),
    .B1(_09718_),
    .B2(_08389_),
    .Y(_09719_));
 sky130_fd_sc_hd__a21oi_4 _15135_ (.A1(_09715_),
    .A2(_09716_),
    .B1(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__o21ai_4 _15136_ (.A1(_09573_),
    .A2(_09711_),
    .B1(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__nor2_2 _15137_ (.A(_08172_),
    .B(net3691),
    .Y(_09722_));
 sky130_fd_sc_hd__o22ai_1 _15138_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .B2(_08171_),
    .Y(_09723_));
 sky130_fd_sc_hd__a211oi_4 _15139_ (.A1(net3949),
    .A2(_09721_),
    .B1(_09722_),
    .C1(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__o21ai_0 _15140_ (.A1(net3626),
    .A2(_09706_),
    .B1(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__xor2_1 _15141_ (.A(_09677_),
    .B(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__nor2_1 _15142_ (.A(net3722),
    .B(_09721_),
    .Y(_09727_));
 sky130_fd_sc_hd__a21oi_1 _15143_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net3722),
    .B1(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_1 _15144_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(net3665),
    .Y(_09729_));
 sky130_fd_sc_hd__o21ai_4 _15145_ (.A1(net3666),
    .A2(_09728_),
    .B1(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__xnor2_1 _15146_ (.A(_08205_),
    .B(_09706_),
    .Y(_09731_));
 sky130_fd_sc_hd__xnor2_1 _15147_ (.A(_09730_),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_1 _15148_ (.A(net3745),
    .B(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__o21ai_4 _15149_ (.A1(net3745),
    .A2(_09726_),
    .B1(_09733_),
    .Y(_09734_));
 sky130_fd_sc_hd__mux2i_1 _15150_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .S(net3928),
    .Y(_09735_));
 sky130_fd_sc_hd__mux2i_1 _15151_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .S(net3928),
    .Y(_09736_));
 sky130_fd_sc_hd__a22oi_1 _15152_ (.A1(net3777),
    .A2(_09735_),
    .B1(_09736_),
    .B2(net3794),
    .Y(_09737_));
 sky130_fd_sc_hd__mux2i_1 _15153_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S(net3928),
    .Y(_09738_));
 sky130_fd_sc_hd__mux2i_1 _15154_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S(net3928),
    .Y(_09739_));
 sky130_fd_sc_hd__a22oi_1 _15155_ (.A1(net3792),
    .A2(_09738_),
    .B1(_09739_),
    .B2(net3779),
    .Y(_09740_));
 sky130_fd_sc_hd__nand3_1 _15156_ (.A(net3774),
    .B(_09737_),
    .C(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__mux4_2 _15157_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net3931),
    .S1(net3911),
    .X(_09742_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net3931),
    .X(_09743_));
 sky130_fd_sc_hd__a221o_1 _15159_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .A2(net320),
    .B1(_09743_),
    .B2(net3911),
    .C1(net3904),
    .X(_09744_));
 sky130_fd_sc_hd__o211ai_1 _15160_ (.A1(_08109_),
    .A2(_09742_),
    .B1(_09744_),
    .C1(net3781),
    .Y(_09745_));
 sky130_fd_sc_hd__mux2i_1 _15161_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .S(net3928),
    .Y(_09746_));
 sky130_fd_sc_hd__mux2i_1 _15162_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S(net3928),
    .Y(_09747_));
 sky130_fd_sc_hd__a22oi_1 _15163_ (.A1(net3777),
    .A2(_09746_),
    .B1(_09747_),
    .B2(net3792),
    .Y(_09748_));
 sky130_fd_sc_hd__mux2i_1 _15164_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .S(net3928),
    .Y(_09749_));
 sky130_fd_sc_hd__mux2i_1 _15165_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S(net3928),
    .Y(_09750_));
 sky130_fd_sc_hd__a22oi_1 _15166_ (.A1(net3794),
    .A2(_09749_),
    .B1(_09750_),
    .B2(net3779),
    .Y(_09751_));
 sky130_fd_sc_hd__nand3_1 _15167_ (.A(_08694_),
    .B(_09748_),
    .C(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__mux2i_1 _15168_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S(net3928),
    .Y(_09753_));
 sky130_fd_sc_hd__mux2i_1 _15169_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .S(net3928),
    .Y(_09754_));
 sky130_fd_sc_hd__a22oi_1 _15170_ (.A1(net3779),
    .A2(_09753_),
    .B1(_09754_),
    .B2(net3794),
    .Y(_09755_));
 sky130_fd_sc_hd__mux2i_1 _15171_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .S(net3928),
    .Y(_09756_));
 sky130_fd_sc_hd__mux2i_1 _15172_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S(net3928),
    .Y(_09757_));
 sky130_fd_sc_hd__a22oi_1 _15173_ (.A1(net3777),
    .A2(_09756_),
    .B1(_09757_),
    .B2(net3792),
    .Y(_09758_));
 sky130_fd_sc_hd__nand3_1 _15174_ (.A(net3784),
    .B(_09755_),
    .C(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__and4_4 _15175_ (.A(_09741_),
    .B(_09745_),
    .C(_09752_),
    .D(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_996 ();
 sky130_fd_sc_hd__o22ai_2 _15178_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .B2(_08171_),
    .Y(_09763_));
 sky130_fd_sc_hd__mux4_2 _15179_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net3894),
    .S1(net303),
    .X(_09764_));
 sky130_fd_sc_hd__nand2_1 _15180_ (.A(net3854),
    .B(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__mux4_2 _15181_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net3894),
    .S1(net303),
    .X(_09766_));
 sky130_fd_sc_hd__nand2_1 _15182_ (.A(_07927_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__and3_4 _15183_ (.A(net3849),
    .B(_09765_),
    .C(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__mux2_1 _15184_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .S(net295),
    .X(_09769_));
 sky130_fd_sc_hd__a22o_1 _15185_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .A2(net3816),
    .B1(_09769_),
    .B2(net3868),
    .X(_09770_));
 sky130_fd_sc_hd__mux2i_1 _15186_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net3868),
    .Y(_09771_));
 sky130_fd_sc_hd__mux2i_1 _15187_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S(net3868),
    .Y(_09772_));
 sky130_fd_sc_hd__o221ai_1 _15188_ (.A1(net362),
    .A2(_09771_),
    .B1(_09772_),
    .B2(_07951_),
    .C1(_07955_),
    .Y(_09773_));
 sky130_fd_sc_hd__a21oi_2 _15189_ (.A1(_07935_),
    .A2(_09770_),
    .B1(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__mux2i_1 _15190_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S(net3878),
    .Y(_09775_));
 sky130_fd_sc_hd__mux2i_1 _15191_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .S(net3878),
    .Y(_09776_));
 sky130_fd_sc_hd__a22oi_1 _15192_ (.A1(net3811),
    .A2(_09775_),
    .B1(_09776_),
    .B2(net3808),
    .Y(_09777_));
 sky130_fd_sc_hd__mux2i_1 _15193_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .S(net3878),
    .Y(_09778_));
 sky130_fd_sc_hd__mux2i_1 _15194_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S(net3878),
    .Y(_09779_));
 sky130_fd_sc_hd__a22oi_1 _15195_ (.A1(net3806),
    .A2(_09778_),
    .B1(_09779_),
    .B2(net3802),
    .Y(_09780_));
 sky130_fd_sc_hd__mux4_2 _15196_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net3894),
    .S1(net3878),
    .X(_09781_));
 sky130_fd_sc_hd__mux4_2 _15197_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net3894),
    .S1(net3878),
    .X(_09782_));
 sky130_fd_sc_hd__a22o_1 _15198_ (.A1(net352),
    .A2(_09781_),
    .B1(_09782_),
    .B2(net3798),
    .X(_09783_));
 sky130_fd_sc_hd__a31oi_2 _15199_ (.A1(net3752),
    .A2(_09777_),
    .A3(_09780_),
    .B1(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__o31ai_4 _15200_ (.A1(net3847),
    .A2(_09774_),
    .A3(_09768_),
    .B1(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__nor2_2 _15201_ (.A(_08172_),
    .B(net3688),
    .Y(_09786_));
 sky130_fd_sc_hd__a211oi_4 _15202_ (.A1(net3949),
    .A2(net3689),
    .B1(_09763_),
    .C1(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__a21oi_4 _15203_ (.A1(net3895),
    .A2(net3700),
    .B1(_09680_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_1 _15204_ (.A(_07888_),
    .B(net3688),
    .Y(_09789_));
 sky130_fd_sc_hd__o21ai_4 _15205_ (.A1(_07888_),
    .A2(_09788_),
    .B1(_09789_),
    .Y(_09790_));
 sky130_fd_sc_hd__nor2_1 _15206_ (.A(net3626),
    .B(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21oi_2 _15207_ (.A1(net3624),
    .A2(_09790_),
    .B1(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__o21a_4 _15208_ (.A1(net3745),
    .A2(_09787_),
    .B1(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__nor2_1 _15209_ (.A(net3722),
    .B(_09760_),
    .Y(_09794_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net3722),
    .B1(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nor2_1 _15211_ (.A(net3666),
    .B(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__a21oi_4 _15212_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(net3665),
    .B1(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__a21oi_2 _15213_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(_07864_),
    .B1(net3745),
    .Y(_09798_));
 sky130_fd_sc_hd__a21oi_4 _15214_ (.A1(net3745),
    .A2(_09797_),
    .B1(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__inv_1 _15215_ (.A(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_2 _15216_ (.A(_09666_),
    .B(_09667_),
    .Y(_09801_));
 sky130_fd_sc_hd__nor2_1 _15217_ (.A(net3755),
    .B(_09593_),
    .Y(_09802_));
 sky130_fd_sc_hd__a21oi_1 _15218_ (.A1(net3755),
    .A2(_09540_),
    .B1(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__nor2_1 _15219_ (.A(net3745),
    .B(_09587_),
    .Y(_09804_));
 sky130_fd_sc_hd__a21oi_1 _15220_ (.A1(net3624),
    .A2(_09566_),
    .B1(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__o21ai_1 _15221_ (.A1(net3626),
    .A2(_09566_),
    .B1(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_2 _15222_ (.A(_09803_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__nor2_1 _15223_ (.A(_09803_),
    .B(_09806_),
    .Y(_09808_));
 sky130_fd_sc_hd__a21oi_1 _15224_ (.A1(_09801_),
    .A2(_09807_),
    .B1(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__a31oi_2 _15225_ (.A1(_09536_),
    .A2(_09597_),
    .A3(_09669_),
    .B1(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__maj3_1 _15226_ (.A(_09793_),
    .B(_09800_),
    .C(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__xor2_2 _15227_ (.A(_09734_),
    .B(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__inv_2 _15228_ (.A(_09812_),
    .Y(net162));
 sky130_fd_sc_hd__xnor2_2 _15229_ (.A(_09793_),
    .B(_09799_),
    .Y(_09813_));
 sky130_fd_sc_hd__xnor2_4 _15230_ (.A(net3511),
    .B(_09813_),
    .Y(net161));
 sky130_fd_sc_hd__nand3_4 _15231_ (.A(_09597_),
    .B(_09734_),
    .C(_09813_),
    .Y(_09814_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_993 ();
 sky130_fd_sc_hd__mux4_2 _15235_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09818_));
 sky130_fd_sc_hd__mux4_2 _15236_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09819_));
 sky130_fd_sc_hd__a22o_4 _15237_ (.A1(_08855_),
    .A2(_09818_),
    .B1(_09819_),
    .B2(_08854_),
    .X(_09820_));
 sky130_fd_sc_hd__mux4_2 _15238_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09821_));
 sky130_fd_sc_hd__nand2_1 _15239_ (.A(net3901),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__mux4_2 _15240_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net3933),
    .S1(net3914),
    .X(_09823_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(_08109_),
    .B(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21oi_2 _15242_ (.A1(_09822_),
    .A2(_09824_),
    .B1(net3768),
    .Y(_09825_));
 sky130_fd_sc_hd__mux2_1 _15243_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .S(net3933),
    .X(_09826_));
 sky130_fd_sc_hd__a221oi_1 _15244_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A2(_08275_),
    .B1(_09826_),
    .B2(net3901),
    .C1(net3914),
    .Y(_09827_));
 sky130_fd_sc_hd__mux4_2 _15245_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net3933),
    .S1(net3901),
    .X(_09828_));
 sky130_fd_sc_hd__o21ai_1 _15246_ (.A1(_08500_),
    .A2(_09828_),
    .B1(net3781),
    .Y(_09829_));
 sky130_fd_sc_hd__mux4_2 _15247_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09830_));
 sky130_fd_sc_hd__mux4_2 _15248_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S0(net3918),
    .S1(net3906),
    .X(_09831_));
 sky130_fd_sc_hd__mux2i_2 _15249_ (.A0(_09830_),
    .A1(_09831_),
    .S(_08109_),
    .Y(_09832_));
 sky130_fd_sc_hd__o22ai_1 _15250_ (.A1(_09827_),
    .A2(_09829_),
    .B1(_09832_),
    .B2(net3769),
    .Y(_09833_));
 sky130_fd_sc_hd__nor3_4 _15251_ (.A(_09833_),
    .B(_09825_),
    .C(_09820_),
    .Y(_09834_));
 sky130_fd_sc_hd__nor2_1 _15252_ (.A(net3722),
    .B(net3687),
    .Y(_09835_));
 sky130_fd_sc_hd__a21oi_1 _15253_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net3722),
    .B1(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__nor2_1 _15254_ (.A(net3666),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__a21oi_4 _15255_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(net3665),
    .B1(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_992 ();
 sky130_fd_sc_hd__a21oi_1 _15257_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_07864_),
    .B1(net3745),
    .Y(_09840_));
 sky130_fd_sc_hd__a21oi_2 _15258_ (.A1(net3745),
    .A2(net436),
    .B1(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__mux4_2 _15259_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net3895),
    .S1(net359),
    .X(_09842_));
 sky130_fd_sc_hd__nand2_1 _15260_ (.A(net3851),
    .B(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__mux4_2 _15261_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net3895),
    .S1(net3858),
    .X(_09844_));
 sky130_fd_sc_hd__nand2_1 _15262_ (.A(_07927_),
    .B(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__and3_4 _15263_ (.A(net3848),
    .B(_09843_),
    .C(_09845_),
    .X(_09846_));
 sky130_fd_sc_hd__mux2_1 _15264_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .S(net3851),
    .X(_09847_));
 sky130_fd_sc_hd__a22o_1 _15265_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A2(net3815),
    .B1(_09847_),
    .B2(net262),
    .X(_09848_));
 sky130_fd_sc_hd__mux2i_1 _15266_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net262),
    .Y(_09849_));
 sky130_fd_sc_hd__mux2i_1 _15267_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S(net262),
    .Y(_09850_));
 sky130_fd_sc_hd__o221ai_1 _15268_ (.A1(net3814),
    .A2(_09849_),
    .B1(_09850_),
    .B2(net429),
    .C1(net3812),
    .Y(_09851_));
 sky130_fd_sc_hd__a21oi_2 _15269_ (.A1(_07935_),
    .A2(_09848_),
    .B1(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__mux2i_1 _15270_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S(net3861),
    .Y(_09853_));
 sky130_fd_sc_hd__mux2i_1 _15271_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .S(net3861),
    .Y(_09854_));
 sky130_fd_sc_hd__a22oi_1 _15272_ (.A1(net3810),
    .A2(_09853_),
    .B1(_09854_),
    .B2(net3809),
    .Y(_09855_));
 sky130_fd_sc_hd__mux2i_1 _15273_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .S(net3861),
    .Y(_09856_));
 sky130_fd_sc_hd__mux2i_1 _15274_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S(net3861),
    .Y(_09857_));
 sky130_fd_sc_hd__a22oi_2 _15275_ (.A1(net3804),
    .A2(_09856_),
    .B1(_09857_),
    .B2(net3803),
    .Y(_09858_));
 sky130_fd_sc_hd__mux4_2 _15276_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net3881),
    .S1(net3861),
    .X(_09859_));
 sky130_fd_sc_hd__mux4_2 _15277_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net3881),
    .S1(net3861),
    .X(_09860_));
 sky130_fd_sc_hd__a22o_4 _15278_ (.A1(net3799),
    .A2(_09859_),
    .B1(_09860_),
    .B2(net3800),
    .X(_09861_));
 sky130_fd_sc_hd__a31oi_4 _15279_ (.A1(net3751),
    .A2(_09855_),
    .A3(_09858_),
    .B1(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__o31ai_4 _15280_ (.A1(net3845),
    .A2(_09846_),
    .A3(_09852_),
    .B1(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__a21oi_2 _15281_ (.A1(net3851),
    .A2(net3700),
    .B1(_09680_),
    .Y(_09864_));
 sky130_fd_sc_hd__nor2_1 _15282_ (.A(net3728),
    .B(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__a21oi_4 _15283_ (.A1(net3728),
    .A2(net3686),
    .B1(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__nor2_1 _15284_ (.A(_08172_),
    .B(net3686),
    .Y(_09867_));
 sky130_fd_sc_hd__o22ai_1 _15285_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .B2(_08171_),
    .Y(_09868_));
 sky130_fd_sc_hd__a211o_1 _15286_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net3687),
    .B1(_09867_),
    .C1(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__a22oi_2 _15287_ (.A1(_08205_),
    .A2(_09866_),
    .B1(_09869_),
    .B2(net3756),
    .Y(_09870_));
 sky130_fd_sc_hd__o21ai_4 _15288_ (.A1(_08442_),
    .A2(_09866_),
    .B1(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__xor2_1 _15289_ (.A(_09841_),
    .B(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__and4b_4 _15290_ (.A_N(_09814_),
    .B(_09872_),
    .C(_09464_),
    .D(_09668_),
    .X(_09873_));
 sky130_fd_sc_hd__maj3_1 _15291_ (.A(_09793_),
    .B(_09800_),
    .C(_09807_),
    .X(_09874_));
 sky130_fd_sc_hd__o22ai_1 _15292_ (.A1(net3626),
    .A2(_09706_),
    .B1(_09724_),
    .B2(net3745),
    .Y(_09875_));
 sky130_fd_sc_hd__a21o_4 _15293_ (.A1(net3624),
    .A2(_09706_),
    .B1(_09875_),
    .X(_09876_));
 sky130_fd_sc_hd__nor2_1 _15294_ (.A(net3755),
    .B(_09730_),
    .Y(_09877_));
 sky130_fd_sc_hd__a21oi_2 _15295_ (.A1(net3755),
    .A2(_09677_),
    .B1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_1 _15296_ (.A(_09876_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__nor2_1 _15297_ (.A(_09876_),
    .B(_09878_),
    .Y(_09880_));
 sky130_fd_sc_hd__a21oi_2 _15298_ (.A1(_09874_),
    .A2(_09879_),
    .B1(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__nor2_1 _15299_ (.A(_09801_),
    .B(_09814_),
    .Y(_09882_));
 sky130_fd_sc_hd__and2_0 _15300_ (.A(_09841_),
    .B(_09871_),
    .X(_09883_));
 sky130_fd_sc_hd__or2_0 _15301_ (.A(_09841_),
    .B(_09871_),
    .X(_09884_));
 sky130_fd_sc_hd__o31a_1 _15302_ (.A1(_09881_),
    .A2(_09882_),
    .A3(_09883_),
    .B1(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__a21oi_4 _15303_ (.A1(_09873_),
    .A2(_09536_),
    .B1(_09885_),
    .Y(_09886_));
 sky130_fd_sc_hd__mux4_2 _15304_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net3926),
    .S1(net3908),
    .X(_09887_));
 sky130_fd_sc_hd__mux4_2 _15305_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net3926),
    .S1(net3908),
    .X(_09888_));
 sky130_fd_sc_hd__mux2_8 _15306_ (.A0(_09887_),
    .A1(_09888_),
    .S(_08109_),
    .X(_09889_));
 sky130_fd_sc_hd__mux2i_1 _15307_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net3931),
    .Y(_09890_));
 sky130_fd_sc_hd__mux2i_1 _15308_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S(net3931),
    .Y(_09891_));
 sky130_fd_sc_hd__a221oi_1 _15309_ (.A1(net3779),
    .A2(_09890_),
    .B1(_09891_),
    .B2(net413),
    .C1(net3899),
    .Y(_09892_));
 sky130_fd_sc_hd__mux2i_1 _15310_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .S(net3931),
    .Y(_09893_));
 sky130_fd_sc_hd__nand3b_1 _15311_ (.A_N(net3904),
    .B(net3932),
    .C(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .Y(_09894_));
 sky130_fd_sc_hd__o211ai_1 _15312_ (.A1(_08109_),
    .A2(_09893_),
    .B1(_09894_),
    .C1(_08500_),
    .Y(_09895_));
 sky130_fd_sc_hd__a221oi_2 _15313_ (.A1(net3899),
    .A2(_09889_),
    .B1(_09892_),
    .B2(_09895_),
    .C1(net3896),
    .Y(_09896_));
 sky130_fd_sc_hd__mux4_2 _15314_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net3928),
    .S1(net3911),
    .X(_09897_));
 sky130_fd_sc_hd__mux4_2 _15315_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net3931),
    .S1(net3911),
    .X(_09898_));
 sky130_fd_sc_hd__o22ai_4 _15316_ (.A1(_09193_),
    .A2(_09897_),
    .B1(_09898_),
    .B2(_09206_),
    .Y(_09899_));
 sky130_fd_sc_hd__mux4_2 _15317_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net3928),
    .S1(net3911),
    .X(_09900_));
 sky130_fd_sc_hd__mux4_2 _15318_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net3928),
    .S1(net3911),
    .X(_09901_));
 sky130_fd_sc_hd__o22ai_4 _15319_ (.A1(_09209_),
    .A2(_09900_),
    .B1(_09901_),
    .B2(_09204_),
    .Y(_09902_));
 sky130_fd_sc_hd__or3_4 _15320_ (.A(_09896_),
    .B(_09899_),
    .C(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__nor2_1 _15321_ (.A(net3722),
    .B(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__a21oi_1 _15322_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net3722),
    .B1(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_2 _15323_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(net3665),
    .Y(_09906_));
 sky130_fd_sc_hd__o21ai_4 _15324_ (.A1(net3666),
    .A2(_09905_),
    .B1(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__nand2_1 _15325_ (.A(net3745),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_990 ();
 sky130_fd_sc_hd__nand3_1 _15328_ (.A(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B(net3739),
    .C(_07864_),
    .Y(_09911_));
 sky130_fd_sc_hd__nand2_2 _15329_ (.A(_09908_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__a21oi_4 _15330_ (.A1(net285),
    .A2(net3700),
    .B1(_09680_),
    .Y(_09913_));
 sky130_fd_sc_hd__mux4_2 _15331_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net3893),
    .S1(net3875),
    .X(_09914_));
 sky130_fd_sc_hd__nand2_1 _15332_ (.A(net3854),
    .B(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__mux4_2 _15333_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net3893),
    .S1(net3875),
    .X(_09916_));
 sky130_fd_sc_hd__nand2_1 _15334_ (.A(_07927_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__and3_4 _15335_ (.A(net3848),
    .B(_09915_),
    .C(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__mux2_1 _15336_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .S(net295),
    .X(_09919_));
 sky130_fd_sc_hd__a22o_1 _15337_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .A2(net345),
    .B1(_09919_),
    .B2(net262),
    .X(_09920_));
 sky130_fd_sc_hd__mux2i_1 _15338_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net262),
    .Y(_09921_));
 sky130_fd_sc_hd__mux2i_1 _15339_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S(net262),
    .Y(_09922_));
 sky130_fd_sc_hd__o22ai_1 _15340_ (.A1(net365),
    .A2(_09921_),
    .B1(_09922_),
    .B2(_07951_),
    .Y(_09923_));
 sky130_fd_sc_hd__a211oi_2 _15341_ (.A1(_07935_),
    .A2(_09920_),
    .B1(_09923_),
    .C1(net3849),
    .Y(_09924_));
 sky130_fd_sc_hd__mux2i_1 _15342_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S(net262),
    .Y(_09925_));
 sky130_fd_sc_hd__mux2i_1 _15343_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .S(net262),
    .Y(_09926_));
 sky130_fd_sc_hd__a22oi_1 _15344_ (.A1(net3811),
    .A2(_09925_),
    .B1(_09926_),
    .B2(net3808),
    .Y(_09927_));
 sky130_fd_sc_hd__mux2i_1 _15345_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .S(net262),
    .Y(_09928_));
 sky130_fd_sc_hd__mux2i_1 _15346_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S(net262),
    .Y(_09929_));
 sky130_fd_sc_hd__a22oi_1 _15347_ (.A1(net3806),
    .A2(_09928_),
    .B1(_09929_),
    .B2(net3802),
    .Y(_09930_));
 sky130_fd_sc_hd__mux4_2 _15348_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net3893),
    .S1(net262),
    .X(_09931_));
 sky130_fd_sc_hd__mux4_2 _15349_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net3893),
    .S1(net262),
    .X(_09932_));
 sky130_fd_sc_hd__a22o_1 _15350_ (.A1(net3798),
    .A2(_09931_),
    .B1(_09932_),
    .B2(net276),
    .X(_09933_));
 sky130_fd_sc_hd__a31oi_2 _15351_ (.A1(net3752),
    .A2(_09927_),
    .A3(_09930_),
    .B1(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__o31ai_4 _15352_ (.A1(net3847),
    .A2(_09918_),
    .A3(_09924_),
    .B1(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_1 _15353_ (.A(net3728),
    .B(net3685),
    .Y(_09936_));
 sky130_fd_sc_hd__o21ai_4 _15354_ (.A1(net3728),
    .A2(_09913_),
    .B1(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__nand2_1 _15355_ (.A(net3624),
    .B(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__nor2_1 _15356_ (.A(_08172_),
    .B(net3685),
    .Y(_09939_));
 sky130_fd_sc_hd__o22ai_1 _15357_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .B2(_08171_),
    .Y(_09940_));
 sky130_fd_sc_hd__a211o_1 _15358_ (.A1(net3949),
    .A2(_09903_),
    .B1(_09939_),
    .C1(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(net3755),
    .B(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__o211ai_1 _15360_ (.A1(net3626),
    .A2(_09937_),
    .B1(_09938_),
    .C1(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__xor2_1 _15361_ (.A(_09912_),
    .B(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__xor2_1 _15362_ (.A(_09886_),
    .B(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__inv_6 _15363_ (.A(net3504),
    .Y(net164));
 sky130_fd_sc_hd__nand3_1 _15364_ (.A(_09314_),
    .B(_09524_),
    .C(_09669_),
    .Y(_09946_));
 sky130_fd_sc_hd__nor2_1 _15365_ (.A(_09814_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__o21ai_0 _15366_ (.A1(net3745),
    .A2(_09787_),
    .B1(_09792_),
    .Y(_09948_));
 sky130_fd_sc_hd__maj3_1 _15367_ (.A(_09665_),
    .B(_09655_),
    .C(_09673_),
    .X(_09949_));
 sky130_fd_sc_hd__nand3_1 _15368_ (.A(_09524_),
    .B(_09537_),
    .C(_09669_),
    .Y(_09950_));
 sky130_fd_sc_hd__a31oi_1 _15369_ (.A1(_09807_),
    .A2(_09949_),
    .A3(_09950_),
    .B1(_09808_),
    .Y(_09951_));
 sky130_fd_sc_hd__maj3_1 _15370_ (.A(_09948_),
    .B(_09799_),
    .C(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__maj3_1 _15371_ (.A(_09876_),
    .B(_09878_),
    .C(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__a31oi_1 _15372_ (.A1(_09376_),
    .A2(_09400_),
    .A3(_09947_),
    .B1(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__xnor2_1 _15373_ (.A(_09872_),
    .B(_09954_),
    .Y(net163));
 sky130_fd_sc_hd__mux2i_1 _15374_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S(net3927),
    .Y(_09955_));
 sky130_fd_sc_hd__mux2i_1 _15375_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .S(net3927),
    .Y(_09956_));
 sky130_fd_sc_hd__a22oi_1 _15376_ (.A1(net3779),
    .A2(_09955_),
    .B1(_09956_),
    .B2(net3794),
    .Y(_09957_));
 sky130_fd_sc_hd__mux2i_1 _15377_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S(net3927),
    .Y(_09958_));
 sky130_fd_sc_hd__mux2i_1 _15378_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .S(net3927),
    .Y(_09959_));
 sky130_fd_sc_hd__a22oi_2 _15379_ (.A1(net3779),
    .A2(_09958_),
    .B1(_09959_),
    .B2(net3794),
    .Y(_09960_));
 sky130_fd_sc_hd__o22ai_4 _15380_ (.A1(_08531_),
    .A2(_09957_),
    .B1(_09960_),
    .B2(_08522_),
    .Y(_09961_));
 sky130_fd_sc_hd__mux2_1 _15381_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S(net3932),
    .X(_09962_));
 sky130_fd_sc_hd__mux2i_1 _15382_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net3932),
    .Y(_09963_));
 sky130_fd_sc_hd__mux2i_1 _15383_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .S(net3932),
    .Y(_09964_));
 sky130_fd_sc_hd__o22ai_1 _15384_ (.A1(net3782),
    .A2(_09963_),
    .B1(_09964_),
    .B2(net3771),
    .Y(_09965_));
 sky130_fd_sc_hd__a21oi_1 _15385_ (.A1(net3792),
    .A2(_09962_),
    .B1(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__a21oi_1 _15386_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A2(net3767),
    .B1(_08538_),
    .Y(_09967_));
 sky130_fd_sc_hd__mux2i_1 _15387_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .S(net3927),
    .Y(_09968_));
 sky130_fd_sc_hd__mux2i_1 _15388_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S(net3927),
    .Y(_09969_));
 sky130_fd_sc_hd__a22oi_1 _15389_ (.A1(net3777),
    .A2(_09968_),
    .B1(_09969_),
    .B2(net3792),
    .Y(_09970_));
 sky130_fd_sc_hd__mux2i_1 _15390_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S(net3927),
    .Y(_09971_));
 sky130_fd_sc_hd__mux2i_1 _15391_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .S(net3927),
    .Y(_09972_));
 sky130_fd_sc_hd__a22oi_1 _15392_ (.A1(net3792),
    .A2(_09971_),
    .B1(_09972_),
    .B2(net3777),
    .Y(_09973_));
 sky130_fd_sc_hd__o22ai_2 _15393_ (.A1(_08531_),
    .A2(_09970_),
    .B1(_09973_),
    .B2(_08522_),
    .Y(_09974_));
 sky130_fd_sc_hd__mux2_1 _15394_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .S(net3928),
    .X(_09975_));
 sky130_fd_sc_hd__mux2i_1 _15395_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S(net3928),
    .Y(_09976_));
 sky130_fd_sc_hd__o21ai_0 _15396_ (.A1(_08261_),
    .A2(_09976_),
    .B1(_08694_),
    .Y(_09977_));
 sky130_fd_sc_hd__mux2i_1 _15397_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .S(net3928),
    .Y(_09978_));
 sky130_fd_sc_hd__mux2i_1 _15398_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .S(net3927),
    .Y(_09979_));
 sky130_fd_sc_hd__o22ai_1 _15399_ (.A1(net3782),
    .A2(_09978_),
    .B1(_09979_),
    .B2(net3771),
    .Y(_09980_));
 sky130_fd_sc_hd__a211oi_1 _15400_ (.A1(net3777),
    .A2(_09975_),
    .B1(_09977_),
    .C1(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__a211o_4 _15401_ (.A1(_09966_),
    .A2(_09967_),
    .B1(_09974_),
    .C1(_09981_),
    .X(_09982_));
 sky130_fd_sc_hd__or2_4 _15402_ (.A(_09961_),
    .B(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__nand2_1 _15403_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .B(net3721),
    .Y(_09984_));
 sky130_fd_sc_hd__o21ai_0 _15404_ (.A1(net3721),
    .A2(_09983_),
    .B1(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__a22o_4 _15405_ (.A1(\cs_registers_i.pc_id_i[24] ),
    .A2(net3665),
    .B1(_09985_),
    .B2(net482),
    .X(_09986_));
 sky130_fd_sc_hd__inv_4 _15406_ (.A(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_989 ();
 sky130_fd_sc_hd__a21oi_1 _15408_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(_07864_),
    .B1(net3745),
    .Y(_09989_));
 sky130_fd_sc_hd__a21oi_2 _15409_ (.A1(net3745),
    .A2(_09987_),
    .B1(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__mux2i_1 _15410_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .S(net3868),
    .Y(_09991_));
 sky130_fd_sc_hd__mux2i_1 _15411_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S(net3868),
    .Y(_09992_));
 sky130_fd_sc_hd__a22oi_1 _15412_ (.A1(net3806),
    .A2(_09991_),
    .B1(_09992_),
    .B2(net3811),
    .Y(_09993_));
 sky130_fd_sc_hd__mux2i_1 _15413_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .S(net3868),
    .Y(_09994_));
 sky130_fd_sc_hd__mux2i_1 _15414_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S(net3868),
    .Y(_09995_));
 sky130_fd_sc_hd__a22oi_1 _15415_ (.A1(net3808),
    .A2(_09994_),
    .B1(_09995_),
    .B2(net3802),
    .Y(_09996_));
 sky130_fd_sc_hd__and3_4 _15416_ (.A(net3752),
    .B(_09993_),
    .C(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__mux2_1 _15417_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net3871),
    .X(_09998_));
 sky130_fd_sc_hd__a221oi_1 _15418_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A2(net3764),
    .B1(_09998_),
    .B2(net322),
    .C1(net3849),
    .Y(_09999_));
 sky130_fd_sc_hd__mux4_2 _15419_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net322),
    .S1(net3868),
    .X(_10000_));
 sky130_fd_sc_hd__nor2_1 _15420_ (.A(_07955_),
    .B(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__nor4_1 _15421_ (.A(net3847),
    .B(net294),
    .C(_09999_),
    .D(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__mux4_2 _15422_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S0(net322),
    .S1(net3868),
    .X(_10003_));
 sky130_fd_sc_hd__mux4_2 _15423_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net322),
    .S1(net3868),
    .X(_10004_));
 sky130_fd_sc_hd__a32oi_1 _15424_ (.A1(net294),
    .A2(_08910_),
    .A3(_10003_),
    .B1(_10004_),
    .B2(net3798),
    .Y(_10005_));
 sky130_fd_sc_hd__mux4_2 _15425_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net322),
    .S1(net262),
    .X(_10006_));
 sky130_fd_sc_hd__mux4_2 _15426_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .S0(net322),
    .S1(net3868),
    .X(_10007_));
 sky130_fd_sc_hd__a32oi_1 _15427_ (.A1(net294),
    .A2(net3765),
    .A3(_10006_),
    .B1(_10007_),
    .B2(net276),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_1 _15428_ (.A(_10005_),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__or3_4 _15429_ (.A(_09997_),
    .B(_10002_),
    .C(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_987 ();
 sky130_fd_sc_hd__o22ai_1 _15432_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .B2(net3786),
    .Y(_10013_));
 sky130_fd_sc_hd__a21oi_1 _15433_ (.A1(net3949),
    .A2(_09983_),
    .B1(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__o21ai_2 _15434_ (.A1(_08172_),
    .A2(_10010_),
    .B1(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__a21oi_2 _15435_ (.A1(net3845),
    .A2(net3700),
    .B1(_09680_),
    .Y(_10016_));
 sky130_fd_sc_hd__nor2_1 _15436_ (.A(net3728),
    .B(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__a21oi_4 _15437_ (.A1(net3728),
    .A2(_10010_),
    .B1(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__nand2_1 _15438_ (.A(_08205_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__o21ai_2 _15439_ (.A1(_08442_),
    .A2(_10018_),
    .B1(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_4 _15440_ (.A1(_07857_),
    .A2(_10015_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__xnor2_2 _15441_ (.A(_09990_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_09944_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__inv_1 _15443_ (.A(_09990_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand2_1 _15444_ (.A(_09912_),
    .B(_09943_),
    .Y(_10025_));
 sky130_fd_sc_hd__maj3_1 _15445_ (.A(_10024_),
    .B(_10021_),
    .C(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__o21ai_2 _15446_ (.A1(_09886_),
    .A2(_10023_),
    .B1(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_986 ();
 sky130_fd_sc_hd__mux2i_1 _15448_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .S(net3870),
    .Y(_10029_));
 sky130_fd_sc_hd__mux2i_1 _15449_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S(net3870),
    .Y(_10030_));
 sky130_fd_sc_hd__a22oi_1 _15450_ (.A1(net3804),
    .A2(_10029_),
    .B1(_10030_),
    .B2(net3811),
    .Y(_10031_));
 sky130_fd_sc_hd__mux2i_1 _15451_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .S(net3870),
    .Y(_10032_));
 sky130_fd_sc_hd__mux2i_1 _15452_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S(net3870),
    .Y(_10033_));
 sky130_fd_sc_hd__a22oi_1 _15453_ (.A1(net3809),
    .A2(_10032_),
    .B1(_10033_),
    .B2(net3803),
    .Y(_10034_));
 sky130_fd_sc_hd__a21oi_1 _15454_ (.A1(_10031_),
    .A2(_10034_),
    .B1(_07955_),
    .Y(_10035_));
 sky130_fd_sc_hd__mux2i_1 _15455_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net3872),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_2 _15456_ (.A(net3813),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__and3_4 _15457_ (.A(net3872),
    .B(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .C(net3804),
    .X(_10038_));
 sky130_fd_sc_hd__mux2i_1 _15458_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S(net3872),
    .Y(_10039_));
 sky130_fd_sc_hd__mux2i_1 _15459_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .S(net3872),
    .Y(_10040_));
 sky130_fd_sc_hd__o22ai_2 _15460_ (.A1(net427),
    .A2(_10039_),
    .B1(_10040_),
    .B2(_08570_),
    .Y(_10041_));
 sky130_fd_sc_hd__o41ai_4 _15461_ (.A1(net3849),
    .A2(_10037_),
    .A3(_10038_),
    .A4(_10041_),
    .B1(_07958_),
    .Y(_10042_));
 sky130_fd_sc_hd__mux4_2 _15462_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .S0(net3872),
    .S1(net294),
    .X(_10043_));
 sky130_fd_sc_hd__mux2i_1 _15463_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S(net3872),
    .Y(_10044_));
 sky130_fd_sc_hd__a21oi_1 _15464_ (.A1(net3803),
    .A2(_10044_),
    .B1(_08650_),
    .Y(_10045_));
 sky130_fd_sc_hd__mux2i_1 _15465_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S(net3870),
    .Y(_10046_));
 sky130_fd_sc_hd__nand2_1 _15466_ (.A(net3811),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__o211ai_1 _15467_ (.A1(net322),
    .A2(_10043_),
    .B1(_10045_),
    .C1(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__mux2i_1 _15468_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .S(net3871),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_2 _15469_ (.A(net3808),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__mux2i_1 _15470_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S(net3871),
    .Y(_10051_));
 sky130_fd_sc_hd__mux2i_1 _15471_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S(net3871),
    .Y(_10052_));
 sky130_fd_sc_hd__a22oi_1 _15472_ (.A1(net3811),
    .A2(_10051_),
    .B1(_10052_),
    .B2(net3803),
    .Y(_10053_));
 sky130_fd_sc_hd__mux2i_1 _15473_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .S(net3871),
    .Y(_10054_));
 sky130_fd_sc_hd__a21oi_2 _15474_ (.A1(net3807),
    .A2(_10054_),
    .B1(_08839_),
    .Y(_10055_));
 sky130_fd_sc_hd__nand3_4 _15475_ (.A(_10050_),
    .B(_10053_),
    .C(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__o211ai_1 _15476_ (.A1(_10035_),
    .A2(_10042_),
    .B1(_10048_),
    .C1(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__a21oi_1 _15477_ (.A1(net3843),
    .A2(net316),
    .B1(_09680_),
    .Y(_10058_));
 sky130_fd_sc_hd__nor2_2 _15478_ (.A(net3728),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__a21oi_4 _15479_ (.A1(net3728),
    .A2(net3684),
    .B1(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__nor2_1 _15480_ (.A(_08442_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__o211a_4 _15481_ (.A1(_10035_),
    .A2(_10042_),
    .B1(_10048_),
    .C1(_10056_),
    .X(_10062_));
 sky130_fd_sc_hd__mux2i_1 _15482_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .S(net267),
    .Y(_10063_));
 sky130_fd_sc_hd__mux2i_1 _15483_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .S(net267),
    .Y(_10064_));
 sky130_fd_sc_hd__a22oi_1 _15484_ (.A1(net3777),
    .A2(_10063_),
    .B1(_10064_),
    .B2(net3793),
    .Y(_10065_));
 sky130_fd_sc_hd__mux2i_1 _15485_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S(net267),
    .Y(_10066_));
 sky130_fd_sc_hd__mux2i_1 _15486_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S(net267),
    .Y(_10067_));
 sky130_fd_sc_hd__a22oi_1 _15487_ (.A1(net3779),
    .A2(_10066_),
    .B1(_10067_),
    .B2(net3792),
    .Y(_10068_));
 sky130_fd_sc_hd__nand3_1 _15488_ (.A(net3773),
    .B(_10065_),
    .C(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__mux4_2 _15489_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net267),
    .S1(net3915),
    .X(_10070_));
 sky130_fd_sc_hd__mux2_1 _15490_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net267),
    .X(_10071_));
 sky130_fd_sc_hd__a221o_1 _15491_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A2(net3788),
    .B1(_10071_),
    .B2(net3915),
    .C1(net3901),
    .X(_10072_));
 sky130_fd_sc_hd__o211ai_1 _15492_ (.A1(_08109_),
    .A2(_10070_),
    .B1(_10072_),
    .C1(net3781),
    .Y(_10073_));
 sky130_fd_sc_hd__mux2i_1 _15493_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .S(net267),
    .Y(_10074_));
 sky130_fd_sc_hd__mux2i_1 _15494_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S(net267),
    .Y(_10075_));
 sky130_fd_sc_hd__a22oi_1 _15495_ (.A1(net3793),
    .A2(_10074_),
    .B1(_10075_),
    .B2(net3779),
    .Y(_10076_));
 sky130_fd_sc_hd__mux2i_1 _15496_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S(net267),
    .Y(_10077_));
 sky130_fd_sc_hd__mux2i_1 _15497_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .S(net267),
    .Y(_10078_));
 sky130_fd_sc_hd__a22oi_1 _15498_ (.A1(net3792),
    .A2(_10077_),
    .B1(_10078_),
    .B2(net3777),
    .Y(_10079_));
 sky130_fd_sc_hd__nand3_1 _15499_ (.A(net3784),
    .B(_10076_),
    .C(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__mux2i_1 _15500_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .S(net3930),
    .Y(_10081_));
 sky130_fd_sc_hd__mux2i_1 _15501_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .S(net3930),
    .Y(_10082_));
 sky130_fd_sc_hd__a22oi_1 _15502_ (.A1(net3777),
    .A2(_10081_),
    .B1(_10082_),
    .B2(net3794),
    .Y(_10083_));
 sky130_fd_sc_hd__mux2i_1 _15503_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S(net3930),
    .Y(_10084_));
 sky130_fd_sc_hd__mux2i_1 _15504_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S(net3930),
    .Y(_10085_));
 sky130_fd_sc_hd__a22oi_1 _15505_ (.A1(net3779),
    .A2(_10084_),
    .B1(_10085_),
    .B2(net3792),
    .Y(_10086_));
 sky130_fd_sc_hd__nand3_2 _15506_ (.A(_08694_),
    .B(_10083_),
    .C(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__and4_4 _15507_ (.A(_10069_),
    .B(_10073_),
    .C(_10080_),
    .D(_10087_),
    .X(_10088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_985 ();
 sky130_fd_sc_hd__o22ai_1 _15509_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .B2(_08171_),
    .Y(_10090_));
 sky130_fd_sc_hd__a221oi_1 _15510_ (.A1(net3736),
    .A2(_10062_),
    .B1(_10088_),
    .B2(net3949),
    .C1(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_08205_),
    .B(_10060_),
    .Y(_10092_));
 sky130_fd_sc_hd__o21ai_2 _15512_ (.A1(net3747),
    .A2(_10091_),
    .B1(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__nor2_4 _15513_ (.A(_10061_),
    .B(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__nor2_1 _15514_ (.A(net3722),
    .B(_10088_),
    .Y(_10095_));
 sky130_fd_sc_hd__a21oi_1 _15515_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net3722),
    .B1(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__nor2_2 _15516_ (.A(net3666),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__a21oi_4 _15517_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(net3665),
    .B1(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nor2_1 _15518_ (.A(net3755),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__a31oi_2 _15519_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net3739),
    .A3(_07864_),
    .B1(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__xnor2_1 _15520_ (.A(_10094_),
    .B(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__xnor2_2 _15521_ (.A(net3502),
    .B(_10101_),
    .Y(net166));
 sky130_fd_sc_hd__nand2_1 _15522_ (.A(_09536_),
    .B(_09669_),
    .Y(_10102_));
 sky130_fd_sc_hd__nor2_1 _15523_ (.A(_09881_),
    .B(_09882_),
    .Y(_10103_));
 sky130_fd_sc_hd__o21ai_0 _15524_ (.A1(_10102_),
    .A2(_09814_),
    .B1(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__maj3_1 _15525_ (.A(_09841_),
    .B(_09871_),
    .C(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__maj3_4 _15526_ (.A(_09912_),
    .B(_09943_),
    .C(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__xor2_4 _15527_ (.A(_10022_),
    .B(_10106_),
    .X(net165));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_984 ();
 sky130_fd_sc_hd__mux4_2 _15529_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net3871),
    .S1(net294),
    .X(_10108_));
 sky130_fd_sc_hd__mux2i_1 _15530_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .S(net294),
    .Y(_10109_));
 sky130_fd_sc_hd__a21oi_1 _15531_ (.A1(net294),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .B1(net3871),
    .Y(_10110_));
 sky130_fd_sc_hd__a211oi_1 _15532_ (.A1(net3871),
    .A2(_10109_),
    .B1(_10110_),
    .C1(net322),
    .Y(_10111_));
 sky130_fd_sc_hd__a21oi_2 _15533_ (.A1(net322),
    .A2(_10108_),
    .B1(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__mux2i_1 _15534_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .S(net3871),
    .Y(_10113_));
 sky130_fd_sc_hd__mux2i_1 _15535_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .S(net3871),
    .Y(_10114_));
 sky130_fd_sc_hd__a22oi_1 _15536_ (.A1(net3806),
    .A2(_10113_),
    .B1(_10114_),
    .B2(net3808),
    .Y(_10115_));
 sky130_fd_sc_hd__mux2i_1 _15537_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S(net3871),
    .Y(_10116_));
 sky130_fd_sc_hd__mux2i_1 _15538_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(net3871),
    .Y(_10117_));
 sky130_fd_sc_hd__a22oi_1 _15539_ (.A1(net3811),
    .A2(_10116_),
    .B1(_10117_),
    .B2(net3802),
    .Y(_10118_));
 sky130_fd_sc_hd__mux4_2 _15540_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net322),
    .S1(net3868),
    .X(_10119_));
 sky130_fd_sc_hd__mux4_2 _15541_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net322),
    .S1(net3868),
    .X(_10120_));
 sky130_fd_sc_hd__a22o_1 _15542_ (.A1(net3798),
    .A2(_10119_),
    .B1(_10120_),
    .B2(net3801),
    .X(_10121_));
 sky130_fd_sc_hd__a31oi_1 _15543_ (.A1(net3765),
    .A2(_10115_),
    .A3(_10118_),
    .B1(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__mux2i_1 _15544_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .S(net3871),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_1 _15545_ (.A(net3808),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__mux2i_1 _15546_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .S(net3871),
    .Y(_10125_));
 sky130_fd_sc_hd__mux2i_1 _15547_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S(net3871),
    .Y(_10126_));
 sky130_fd_sc_hd__a22oi_1 _15548_ (.A1(net3806),
    .A2(_10125_),
    .B1(_10126_),
    .B2(net3811),
    .Y(_10127_));
 sky130_fd_sc_hd__mux2i_1 _15549_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S(net3871),
    .Y(_10128_));
 sky130_fd_sc_hd__a21oi_1 _15550_ (.A1(net3803),
    .A2(_10128_),
    .B1(_08650_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand3_1 _15551_ (.A(_10124_),
    .B(_10127_),
    .C(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__o211ai_1 _15552_ (.A1(_09038_),
    .A2(_10112_),
    .B1(_10122_),
    .C1(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__mux2i_1 _15553_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .S(net3930),
    .Y(_10132_));
 sky130_fd_sc_hd__mux2i_1 _15554_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .S(net3930),
    .Y(_10133_));
 sky130_fd_sc_hd__a22oi_1 _15555_ (.A1(net3777),
    .A2(_10132_),
    .B1(_10133_),
    .B2(net3794),
    .Y(_10134_));
 sky130_fd_sc_hd__mux2i_1 _15556_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S(net3930),
    .Y(_10135_));
 sky130_fd_sc_hd__mux2i_1 _15557_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S(net3930),
    .Y(_10136_));
 sky130_fd_sc_hd__a22oi_1 _15558_ (.A1(net3779),
    .A2(_10135_),
    .B1(_10136_),
    .B2(net3792),
    .Y(_10137_));
 sky130_fd_sc_hd__nand3_1 _15559_ (.A(_08694_),
    .B(_10134_),
    .C(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__mux4_2 _15560_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net267),
    .S1(net3914),
    .X(_10139_));
 sky130_fd_sc_hd__mux2_1 _15561_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net267),
    .X(_10140_));
 sky130_fd_sc_hd__a221o_1 _15562_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .A2(net3788),
    .B1(_10140_),
    .B2(net3914),
    .C1(net3904),
    .X(_10141_));
 sky130_fd_sc_hd__o211ai_1 _15563_ (.A1(_08109_),
    .A2(_10139_),
    .B1(_10141_),
    .C1(net3781),
    .Y(_10142_));
 sky130_fd_sc_hd__mux2i_1 _15564_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .S(net3930),
    .Y(_10143_));
 sky130_fd_sc_hd__mux2i_1 _15565_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .S(net3930),
    .Y(_10144_));
 sky130_fd_sc_hd__a22oi_1 _15566_ (.A1(net3794),
    .A2(_10143_),
    .B1(_10144_),
    .B2(net3777),
    .Y(_10145_));
 sky130_fd_sc_hd__mux2i_1 _15567_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S(net3930),
    .Y(_10146_));
 sky130_fd_sc_hd__mux2i_1 _15568_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S(net3930),
    .Y(_10147_));
 sky130_fd_sc_hd__a22oi_1 _15569_ (.A1(net3792),
    .A2(_10146_),
    .B1(_10147_),
    .B2(net3779),
    .Y(_10148_));
 sky130_fd_sc_hd__nand3_1 _15570_ (.A(net3773),
    .B(_10145_),
    .C(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__mux2i_1 _15571_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .S(net3930),
    .Y(_10150_));
 sky130_fd_sc_hd__mux2i_1 _15572_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S(net3930),
    .Y(_10151_));
 sky130_fd_sc_hd__a22oi_1 _15573_ (.A1(net3794),
    .A2(_10150_),
    .B1(_10151_),
    .B2(net3779),
    .Y(_10152_));
 sky130_fd_sc_hd__mux2i_1 _15574_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(net3930),
    .Y(_10153_));
 sky130_fd_sc_hd__mux2i_1 _15575_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .S(net3930),
    .Y(_10154_));
 sky130_fd_sc_hd__a22oi_1 _15576_ (.A1(net3792),
    .A2(_10153_),
    .B1(_10154_),
    .B2(net3777),
    .Y(_10155_));
 sky130_fd_sc_hd__nand3_1 _15577_ (.A(net3784),
    .B(_10152_),
    .C(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__and4_4 _15578_ (.A(_10138_),
    .B(_10142_),
    .C(_10149_),
    .D(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_982 ();
 sky130_fd_sc_hd__o22ai_1 _15581_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .B2(_08171_),
    .Y(_10160_));
 sky130_fd_sc_hd__a21oi_1 _15582_ (.A1(net3949),
    .A2(net3682),
    .B1(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__o21ai_2 _15583_ (.A1(_08172_),
    .A2(net3683),
    .B1(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__a21oi_1 _15584_ (.A1(net3842),
    .A2(net316),
    .B1(_09680_),
    .Y(_10163_));
 sky130_fd_sc_hd__nor2_1 _15585_ (.A(_07888_),
    .B(_10163_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21oi_4 _15586_ (.A1(_07888_),
    .A2(net3683),
    .B1(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__nand2_1 _15587_ (.A(_08205_),
    .B(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__o21ai_2 _15588_ (.A1(_08442_),
    .A2(_10165_),
    .B1(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__a21oi_4 _15589_ (.A1(_07857_),
    .A2(_10162_),
    .B1(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_981 ();
 sky130_fd_sc_hd__nor2_1 _15591_ (.A(net3721),
    .B(_10157_),
    .Y(_10170_));
 sky130_fd_sc_hd__a21oi_1 _15592_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net3721),
    .B1(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__nor2_2 _15593_ (.A(net3666),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__a21oi_4 _15594_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(net3665),
    .B1(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor2_1 _15595_ (.A(net3755),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__a31oi_2 _15596_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net3739),
    .A3(_07864_),
    .B1(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__o22ai_2 _15597_ (.A1(_10094_),
    .A2(_10100_),
    .B1(_10168_),
    .B2(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_1 _15598_ (.A(_10094_),
    .B(_10100_),
    .Y(_10177_));
 sky130_fd_sc_hd__nand2_1 _15599_ (.A(_10168_),
    .B(_10175_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_1 _15600_ (.A(_10177_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__o21ai_1 _15601_ (.A1(_10168_),
    .A2(_10175_),
    .B1(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__o21ai_2 _15602_ (.A1(net3502),
    .A2(_10176_),
    .B1(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_979 ();
 sky130_fd_sc_hd__mux4_2 _15605_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net3931),
    .S1(net3911),
    .X(_10184_));
 sky130_fd_sc_hd__mux4_2 _15606_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net3927),
    .S1(net3911),
    .X(_10185_));
 sky130_fd_sc_hd__o22ai_1 _15607_ (.A1(_09193_),
    .A2(_10184_),
    .B1(_10185_),
    .B2(_09206_),
    .Y(_10186_));
 sky130_fd_sc_hd__mux4_2 _15608_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net3928),
    .S1(net3911),
    .X(_10187_));
 sky130_fd_sc_hd__mux4_2 _15609_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net3928),
    .S1(net3911),
    .X(_10188_));
 sky130_fd_sc_hd__o22ai_1 _15610_ (.A1(_09209_),
    .A2(_10187_),
    .B1(_10188_),
    .B2(_09204_),
    .Y(_10189_));
 sky130_fd_sc_hd__mux2i_1 _15611_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .S(net3932),
    .Y(_10190_));
 sky130_fd_sc_hd__mux2i_1 _15612_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S(net3932),
    .Y(_10191_));
 sky130_fd_sc_hd__o22ai_1 _15613_ (.A1(net3771),
    .A2(_10190_),
    .B1(_10191_),
    .B2(net3783),
    .Y(_10192_));
 sky130_fd_sc_hd__mux2i_1 _15614_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net3932),
    .Y(_10193_));
 sky130_fd_sc_hd__o2bb2ai_1 _15615_ (.A1_N(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .A2_N(net3767),
    .B1(_10193_),
    .B2(net3782),
    .Y(_10194_));
 sky130_fd_sc_hd__nor3_1 _15616_ (.A(_08538_),
    .B(_10192_),
    .C(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__mux4_2 _15617_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net3927),
    .S1(net3911),
    .X(_10196_));
 sky130_fd_sc_hd__mux4_2 _15618_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net3927),
    .S1(net3911),
    .X(_10197_));
 sky130_fd_sc_hd__o22ai_2 _15619_ (.A1(net3770),
    .A2(_10196_),
    .B1(_10197_),
    .B2(_08389_),
    .Y(_10198_));
 sky130_fd_sc_hd__or4_4 _15620_ (.A(_10186_),
    .B(_10189_),
    .C(_10195_),
    .D(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__nor2_1 _15621_ (.A(net3723),
    .B(net3681),
    .Y(_10200_));
 sky130_fd_sc_hd__a21oi_1 _15622_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net3723),
    .B1(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_2 _15623_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(net3665),
    .Y(_10202_));
 sky130_fd_sc_hd__o21ai_4 _15624_ (.A1(net269),
    .A2(_10201_),
    .B1(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__inv_6 _15625_ (.A(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .Y(_10204_));
 sky130_fd_sc_hd__nor3_4 _15626_ (.A(_10204_),
    .B(net3747),
    .C(net3786),
    .Y(_10205_));
 sky130_fd_sc_hd__a21oi_2 _15627_ (.A1(net3745),
    .A2(_10203_),
    .B1(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__mux2_1 _15628_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net3868),
    .X(_10207_));
 sky130_fd_sc_hd__a221oi_1 _15629_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .A2(net3764),
    .B1(_10207_),
    .B2(net322),
    .C1(net294),
    .Y(_10208_));
 sky130_fd_sc_hd__mux4_2 _15630_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net322),
    .S1(net3868),
    .X(_10209_));
 sky130_fd_sc_hd__o21ai_0 _15631_ (.A1(_07927_),
    .A2(_10209_),
    .B1(net3762),
    .Y(_10210_));
 sky130_fd_sc_hd__mux4_2 _15632_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net3893),
    .S1(net3879),
    .X(_10211_));
 sky130_fd_sc_hd__mux4_2 _15633_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net3893),
    .S1(net262),
    .X(_10212_));
 sky130_fd_sc_hd__a32oi_1 _15634_ (.A1(net294),
    .A2(net3765),
    .A3(_10211_),
    .B1(_10212_),
    .B2(net3798),
    .Y(_10213_));
 sky130_fd_sc_hd__o21ai_2 _15635_ (.A1(_10208_),
    .A2(_10210_),
    .B1(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__nor2_4 _15636_ (.A(net3844),
    .B(net322),
    .Y(_10215_));
 sky130_fd_sc_hd__mux2i_2 _15637_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .S(net3877),
    .Y(_10216_));
 sky130_fd_sc_hd__mux2i_1 _15638_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .S(net3877),
    .Y(_10217_));
 sky130_fd_sc_hd__mux4_2 _15639_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net3877),
    .S1(net3847),
    .X(_10218_));
 sky130_fd_sc_hd__o2bb2ai_2 _15640_ (.A1_N(net3763),
    .A2_N(_10217_),
    .B1(_10218_),
    .B2(_07935_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand2b_4 _15641_ (.A_N(net3854),
    .B(net3848),
    .Y(_10220_));
 sky130_fd_sc_hd__a211oi_4 _15642_ (.A1(_10215_),
    .A2(_10216_),
    .B1(_10219_),
    .C1(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__mux2i_1 _15643_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .S(net262),
    .Y(_10222_));
 sky130_fd_sc_hd__mux2i_1 _15644_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S(net262),
    .Y(_10223_));
 sky130_fd_sc_hd__a22oi_1 _15645_ (.A1(net3806),
    .A2(_10222_),
    .B1(_10223_),
    .B2(net3811),
    .Y(_10224_));
 sky130_fd_sc_hd__mux2i_1 _15646_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .S(net262),
    .Y(_10225_));
 sky130_fd_sc_hd__mux2i_1 _15647_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S(net262),
    .Y(_10226_));
 sky130_fd_sc_hd__a22oi_1 _15648_ (.A1(net3808),
    .A2(_10225_),
    .B1(_10226_),
    .B2(net3802),
    .Y(_10227_));
 sky130_fd_sc_hd__nand3_2 _15649_ (.A(net3752),
    .B(_10224_),
    .C(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__nor3b_4 _15650_ (.A(_10214_),
    .B(_10221_),
    .C_N(_10228_),
    .Y(_10229_));
 sky130_fd_sc_hd__a211oi_2 _15651_ (.A1(net3841),
    .A2(net316),
    .B1(_09680_),
    .C1(net3728),
    .Y(_10230_));
 sky130_fd_sc_hd__a21oi_4 _15652_ (.A1(_07888_),
    .A2(net3680),
    .B1(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_978 ();
 sky130_fd_sc_hd__o22ai_1 _15654_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .B2(net3786),
    .Y(_10233_));
 sky130_fd_sc_hd__a221oi_1 _15655_ (.A1(net3949),
    .A2(net3681),
    .B1(net3680),
    .B2(net3736),
    .C1(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__o22ai_2 _15656_ (.A1(net3626),
    .A2(_10231_),
    .B1(_10234_),
    .B2(net3747),
    .Y(_10235_));
 sky130_fd_sc_hd__a21oi_4 _15657_ (.A1(net3624),
    .A2(_10231_),
    .B1(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__xor2_1 _15658_ (.A(_10206_),
    .B(_10236_),
    .X(_10237_));
 sky130_fd_sc_hd__xor2_2 _15659_ (.A(_10181_),
    .B(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__inv_6 _15660_ (.A(_10238_),
    .Y(net168));
 sky130_fd_sc_hd__xnor2_1 _15661_ (.A(_10168_),
    .B(_10175_),
    .Y(_10239_));
 sky130_fd_sc_hd__nor2_1 _15662_ (.A(_10094_),
    .B(_10100_),
    .Y(_10240_));
 sky130_fd_sc_hd__o21ai_0 _15663_ (.A1(net3502),
    .A2(_10240_),
    .B1(_10177_),
    .Y(_10241_));
 sky130_fd_sc_hd__xnor2_1 _15664_ (.A(_10239_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__inv_2 _15665_ (.A(net323),
    .Y(net167));
 sky130_fd_sc_hd__mux2i_1 _15666_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .S(net3924),
    .Y(_10243_));
 sky130_fd_sc_hd__mux2i_1 _15667_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .S(net3924),
    .Y(_10244_));
 sky130_fd_sc_hd__a22oi_1 _15668_ (.A1(net3776),
    .A2(_10243_),
    .B1(_10244_),
    .B2(net3795),
    .Y(_10245_));
 sky130_fd_sc_hd__mux2i_1 _15669_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S(net3924),
    .Y(_10246_));
 sky130_fd_sc_hd__mux2i_1 _15670_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S(net3924),
    .Y(_10247_));
 sky130_fd_sc_hd__a22oi_1 _15671_ (.A1(net3778),
    .A2(_10246_),
    .B1(_10247_),
    .B2(net3790),
    .Y(_10248_));
 sky130_fd_sc_hd__and3_1 _15672_ (.A(net3784),
    .B(_10245_),
    .C(_10248_),
    .X(_10249_));
 sky130_fd_sc_hd__mux2i_1 _15673_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S(net3921),
    .Y(_10250_));
 sky130_fd_sc_hd__mux2i_1 _15674_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .S(net3921),
    .Y(_10251_));
 sky130_fd_sc_hd__a22oi_1 _15675_ (.A1(net3778),
    .A2(_10250_),
    .B1(_10251_),
    .B2(net3795),
    .Y(_10252_));
 sky130_fd_sc_hd__mux2i_1 _15676_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .S(net3921),
    .Y(_10253_));
 sky130_fd_sc_hd__mux2i_1 _15677_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S(net3921),
    .Y(_10254_));
 sky130_fd_sc_hd__a22oi_1 _15678_ (.A1(net3776),
    .A2(_10253_),
    .B1(_10254_),
    .B2(net3790),
    .Y(_10255_));
 sky130_fd_sc_hd__and3_4 _15679_ (.A(net3774),
    .B(_10252_),
    .C(_10255_),
    .X(_10256_));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net3923),
    .X(_10257_));
 sky130_fd_sc_hd__a221oi_1 _15681_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A2(net319),
    .B1(_10257_),
    .B2(net3910),
    .C1(net3905),
    .Y(_10258_));
 sky130_fd_sc_hd__mux4_2 _15682_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net3923),
    .S1(net3910),
    .X(_10259_));
 sky130_fd_sc_hd__o21ai_0 _15683_ (.A1(_08109_),
    .A2(_10259_),
    .B1(net3781),
    .Y(_10260_));
 sky130_fd_sc_hd__mux4_2 _15684_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net3920),
    .S1(net3907),
    .X(_10261_));
 sky130_fd_sc_hd__mux4_2 _15685_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net3920),
    .S1(net3907),
    .X(_10262_));
 sky130_fd_sc_hd__a22oi_2 _15686_ (.A1(_08855_),
    .A2(_10261_),
    .B1(_10262_),
    .B2(_08854_),
    .Y(_10263_));
 sky130_fd_sc_hd__o21ai_2 _15687_ (.A1(_10258_),
    .A2(_10260_),
    .B1(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__nor3_2 _15688_ (.A(_10249_),
    .B(_10256_),
    .C(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(net3723),
    .B(net3678),
    .Y(_10266_));
 sky130_fd_sc_hd__a21oi_1 _15690_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net3723),
    .B1(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__nor2_2 _15691_ (.A(net269),
    .B(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__a21oi_4 _15692_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(net3665),
    .B1(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_977 ();
 sky130_fd_sc_hd__a21oi_1 _15694_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(_07864_),
    .B1(net3745),
    .Y(_10271_));
 sky130_fd_sc_hd__a21oi_2 _15695_ (.A1(net3745),
    .A2(_10269_),
    .B1(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__mux2_1 _15696_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net3865),
    .X(_10273_));
 sky130_fd_sc_hd__a221oi_1 _15697_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A2(net3764),
    .B1(_10273_),
    .B2(net3889),
    .C1(net3855),
    .Y(_10274_));
 sky130_fd_sc_hd__mux4_2 _15698_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net3889),
    .S1(net3865),
    .X(_10275_));
 sky130_fd_sc_hd__nor2_1 _15699_ (.A(_07927_),
    .B(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__mux2i_1 _15700_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S(net3863),
    .Y(_10277_));
 sky130_fd_sc_hd__mux2i_1 _15701_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .S(net3863),
    .Y(_10278_));
 sky130_fd_sc_hd__a22oi_1 _15702_ (.A1(net3811),
    .A2(_10277_),
    .B1(_10278_),
    .B2(net3808),
    .Y(_10279_));
 sky130_fd_sc_hd__mux2i_1 _15703_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .S(net3863),
    .Y(_10280_));
 sky130_fd_sc_hd__mux2i_1 _15704_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S(net3863),
    .Y(_10281_));
 sky130_fd_sc_hd__a22oi_1 _15705_ (.A1(net3805),
    .A2(_10280_),
    .B1(_10281_),
    .B2(net3802),
    .Y(_10282_));
 sky130_fd_sc_hd__mux4_2 _15706_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net3883),
    .S1(net3863),
    .X(_10283_));
 sky130_fd_sc_hd__mux4_2 _15707_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net3883),
    .S1(net3863),
    .X(_10284_));
 sky130_fd_sc_hd__a22o_4 _15708_ (.A1(net3800),
    .A2(_10283_),
    .B1(_10284_),
    .B2(net3799),
    .X(_10285_));
 sky130_fd_sc_hd__a31oi_2 _15709_ (.A1(net3752),
    .A2(_10279_),
    .A3(_10282_),
    .B1(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__mux2i_1 _15710_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .S(net3863),
    .Y(_10287_));
 sky130_fd_sc_hd__mux2i_1 _15711_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S(net3863),
    .Y(_10288_));
 sky130_fd_sc_hd__a22oi_1 _15712_ (.A1(net3805),
    .A2(_10287_),
    .B1(_10288_),
    .B2(net3811),
    .Y(_10289_));
 sky130_fd_sc_hd__mux2i_1 _15713_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .S(net3863),
    .Y(_10290_));
 sky130_fd_sc_hd__mux2i_1 _15714_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S(net3863),
    .Y(_10291_));
 sky130_fd_sc_hd__a22oi_1 _15715_ (.A1(net3808),
    .A2(_10290_),
    .B1(_10291_),
    .B2(net3802),
    .Y(_10292_));
 sky130_fd_sc_hd__nand3_1 _15716_ (.A(net3766),
    .B(_10289_),
    .C(_10292_),
    .Y(_10293_));
 sky130_fd_sc_hd__o311a_4 _15717_ (.A1(_09038_),
    .A2(_10274_),
    .A3(_10276_),
    .B1(_10286_),
    .C1(_10293_),
    .X(_10294_));
 sky130_fd_sc_hd__a211oi_1 _15718_ (.A1(net3840),
    .A2(net316),
    .B1(_09680_),
    .C1(net3728),
    .Y(_10295_));
 sky130_fd_sc_hd__a21o_4 _15719_ (.A1(net3728),
    .A2(_10294_),
    .B1(_10295_),
    .X(_10296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_976 ();
 sky130_fd_sc_hd__o22ai_1 _15721_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .B2(net3786),
    .Y(_10298_));
 sky130_fd_sc_hd__a221oi_1 _15722_ (.A1(net3949),
    .A2(net3679),
    .B1(_10294_),
    .B2(net3736),
    .C1(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__nor2_2 _15723_ (.A(net3747),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__a21oi_1 _15724_ (.A1(_08205_),
    .A2(_10296_),
    .B1(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_4 _15725_ (.A1(_08442_),
    .A2(_10296_),
    .B1(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__nor2_1 _15726_ (.A(_10206_),
    .B(_10236_),
    .Y(_10303_));
 sky130_fd_sc_hd__nand2_1 _15727_ (.A(_10206_),
    .B(_10236_),
    .Y(_10304_));
 sky130_fd_sc_hd__a21oi_1 _15728_ (.A1(_10180_),
    .A2(_10304_),
    .B1(_10303_),
    .Y(_10305_));
 sky130_fd_sc_hd__inv_1 _15729_ (.A(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__o31a_4 _15730_ (.A1(_10303_),
    .A2(_10176_),
    .A3(_10027_),
    .B1(_10306_),
    .X(_10307_));
 sky130_fd_sc_hd__maj3_4 _15731_ (.A(_10272_),
    .B(_10302_),
    .C(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_975 ();
 sky130_fd_sc_hd__mux2i_1 _15733_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .S(net267),
    .Y(_10310_));
 sky130_fd_sc_hd__mux2i_1 _15734_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S(net267),
    .Y(_10311_));
 sky130_fd_sc_hd__a22oi_1 _15735_ (.A1(net260),
    .A2(_10310_),
    .B1(_10311_),
    .B2(net3791),
    .Y(_10312_));
 sky130_fd_sc_hd__mux2i_1 _15736_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .S(net267),
    .Y(_10313_));
 sky130_fd_sc_hd__mux2i_1 _15737_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S(net267),
    .Y(_10314_));
 sky130_fd_sc_hd__a22oi_1 _15738_ (.A1(net3793),
    .A2(_10313_),
    .B1(_10314_),
    .B2(net3780),
    .Y(_10315_));
 sky130_fd_sc_hd__and3_4 _15739_ (.A(net3784),
    .B(_10312_),
    .C(_10315_),
    .X(_10316_));
 sky130_fd_sc_hd__mux2i_1 _15740_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S(net3919),
    .Y(_10317_));
 sky130_fd_sc_hd__mux2i_1 _15741_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .S(net3919),
    .Y(_10318_));
 sky130_fd_sc_hd__a22oi_1 _15742_ (.A1(net3780),
    .A2(_10317_),
    .B1(_10318_),
    .B2(net3793),
    .Y(_10319_));
 sky130_fd_sc_hd__mux2i_1 _15743_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .S(net3919),
    .Y(_10320_));
 sky130_fd_sc_hd__mux2i_1 _15744_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(net346),
    .Y(_10321_));
 sky130_fd_sc_hd__a22oi_1 _15745_ (.A1(net260),
    .A2(_10320_),
    .B1(_10321_),
    .B2(net411),
    .Y(_10322_));
 sky130_fd_sc_hd__and3_4 _15746_ (.A(net3773),
    .B(_10319_),
    .C(_10322_),
    .X(_10323_));
 sky130_fd_sc_hd__mux2_1 _15747_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net267),
    .X(_10324_));
 sky130_fd_sc_hd__a221oi_1 _15748_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A2(net3789),
    .B1(_10324_),
    .B2(net3914),
    .C1(net3901),
    .Y(_10325_));
 sky130_fd_sc_hd__mux4_2 _15749_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net3933),
    .S1(net3914),
    .X(_10326_));
 sky130_fd_sc_hd__o21ai_2 _15750_ (.A1(_08109_),
    .A2(_10326_),
    .B1(net3781),
    .Y(_10327_));
 sky130_fd_sc_hd__mux4_2 _15751_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net3918),
    .S1(net3908),
    .X(_10328_));
 sky130_fd_sc_hd__mux4_2 _15752_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net3919),
    .S1(net3908),
    .X(_10329_));
 sky130_fd_sc_hd__a22oi_1 _15753_ (.A1(_08855_),
    .A2(_10328_),
    .B1(_10329_),
    .B2(_08854_),
    .Y(_10330_));
 sky130_fd_sc_hd__o21ai_2 _15754_ (.A1(_10325_),
    .A2(_10327_),
    .B1(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__nor3_4 _15755_ (.A(_10316_),
    .B(_10323_),
    .C(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__nor2_1 _15756_ (.A(net3722),
    .B(net3676),
    .Y(_10333_));
 sky130_fd_sc_hd__a21oi_1 _15757_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net3722),
    .B1(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__nor2_2 _15758_ (.A(net3666),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__a21oi_4 _15759_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(net3665),
    .B1(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__nor2_1 _15760_ (.A(net3755),
    .B(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__a31oi_2 _15761_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net3739),
    .A3(_07864_),
    .B1(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__mux2i_1 _15762_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .S(net3861),
    .Y(_10339_));
 sky130_fd_sc_hd__mux2i_1 _15763_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S(net3861),
    .Y(_10340_));
 sky130_fd_sc_hd__a22oi_1 _15764_ (.A1(net3804),
    .A2(_10339_),
    .B1(_10340_),
    .B2(net3810),
    .Y(_10341_));
 sky130_fd_sc_hd__mux2i_1 _15765_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .S(net3861),
    .Y(_10342_));
 sky130_fd_sc_hd__mux2i_1 _15766_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(net3861),
    .Y(_10343_));
 sky130_fd_sc_hd__a22oi_1 _15767_ (.A1(net3809),
    .A2(_10342_),
    .B1(_10343_),
    .B2(net3803),
    .Y(_10344_));
 sky130_fd_sc_hd__and3_4 _15768_ (.A(net3751),
    .B(_10341_),
    .C(_10344_),
    .X(_10345_));
 sky130_fd_sc_hd__mux2_1 _15769_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net3866),
    .X(_10346_));
 sky130_fd_sc_hd__a221oi_1 _15770_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A2(net3764),
    .B1(_10346_),
    .B2(net322),
    .C1(net294),
    .Y(_10347_));
 sky130_fd_sc_hd__mux4_2 _15771_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net3895),
    .S1(net359),
    .X(_10348_));
 sky130_fd_sc_hd__o21ai_0 _15772_ (.A1(_07927_),
    .A2(_10348_),
    .B1(net3762),
    .Y(_10349_));
 sky130_fd_sc_hd__mux4_2 _15773_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net322),
    .S1(net3861),
    .X(_10350_));
 sky130_fd_sc_hd__mux4_2 _15774_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net3882),
    .S1(net3861),
    .X(_10351_));
 sky130_fd_sc_hd__a32oi_2 _15775_ (.A1(net3852),
    .A2(net3766),
    .A3(_10350_),
    .B1(_10351_),
    .B2(net3799),
    .Y(_10352_));
 sky130_fd_sc_hd__o21ai_2 _15776_ (.A1(_10347_),
    .A2(_10349_),
    .B1(_10352_),
    .Y(_10353_));
 sky130_fd_sc_hd__mux4_2 _15777_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net3861),
    .S1(net3845),
    .X(_10354_));
 sky130_fd_sc_hd__mux2i_1 _15778_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .S(net3866),
    .Y(_10355_));
 sky130_fd_sc_hd__a21oi_1 _15779_ (.A1(_10215_),
    .A2(_10355_),
    .B1(_10220_),
    .Y(_10356_));
 sky130_fd_sc_hd__mux2i_1 _15780_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .S(net3861),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_1 _15781_ (.A(net3763),
    .B(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__o211ai_1 _15782_ (.A1(_07935_),
    .A2(_10354_),
    .B1(_10356_),
    .C1(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__or3b_4 _15783_ (.A(_10345_),
    .B(_10353_),
    .C_N(_10359_),
    .X(_10360_));
 sky130_fd_sc_hd__o22ai_1 _15784_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .B2(_08171_),
    .Y(_10361_));
 sky130_fd_sc_hd__a21oi_1 _15785_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net3676),
    .B1(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__o21ai_2 _15786_ (.A1(_08172_),
    .A2(_10360_),
    .B1(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__a21oi_1 _15787_ (.A1(net3839),
    .A2(net316),
    .B1(_09680_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_2 _15788_ (.A(net3718),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__o21ai_4 _15789_ (.A1(net3718),
    .A2(_10360_),
    .B1(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_1 _15790_ (.A(_08205_),
    .B(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__o21ai_2 _15791_ (.A1(_08442_),
    .A2(_10366_),
    .B1(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__a21oi_4 _15792_ (.A1(net3756),
    .A2(_10363_),
    .B1(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__xnor2_1 _15793_ (.A(_10338_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__xnor2_4 _15794_ (.A(_10308_),
    .B(_10370_),
    .Y(net170));
 sky130_fd_sc_hd__xor2_1 _15795_ (.A(_10272_),
    .B(_10302_),
    .X(_10371_));
 sky130_fd_sc_hd__xnor2_4 _15796_ (.A(net468),
    .B(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__inv_16 _15797_ (.A(_10372_),
    .Y(net169));
 sky130_fd_sc_hd__mux4_2 _15798_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .S0(net3885),
    .S1(net294),
    .X(_10373_));
 sky130_fd_sc_hd__mux4_2 _15799_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S0(net3885),
    .S1(net294),
    .X(_10374_));
 sky130_fd_sc_hd__mux2i_1 _15800_ (.A0(_10373_),
    .A1(_10374_),
    .S(net262),
    .Y(_10375_));
 sky130_fd_sc_hd__mux2i_1 _15801_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .S(net3870),
    .Y(_10376_));
 sky130_fd_sc_hd__mux2i_1 _15802_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S(net3870),
    .Y(_10377_));
 sky130_fd_sc_hd__a22oi_1 _15803_ (.A1(net3809),
    .A2(_10376_),
    .B1(_10377_),
    .B2(net3810),
    .Y(_10378_));
 sky130_fd_sc_hd__mux2i_1 _15804_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .S(net3870),
    .Y(_10379_));
 sky130_fd_sc_hd__mux2i_1 _15805_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S(net3871),
    .Y(_10380_));
 sky130_fd_sc_hd__a22oi_1 _15806_ (.A1(net3804),
    .A2(_10379_),
    .B1(_10380_),
    .B2(net3803),
    .Y(_10381_));
 sky130_fd_sc_hd__mux4_2 _15807_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net3885),
    .S1(net262),
    .X(_10382_));
 sky130_fd_sc_hd__mux4_2 _15808_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net3885),
    .S1(net262),
    .X(_10383_));
 sky130_fd_sc_hd__a22o_1 _15809_ (.A1(net3798),
    .A2(_10382_),
    .B1(_10383_),
    .B2(net3801),
    .X(_10384_));
 sky130_fd_sc_hd__a31oi_1 _15810_ (.A1(net3751),
    .A2(_10378_),
    .A3(_10381_),
    .B1(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__mux4_2 _15811_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net3885),
    .S1(net262),
    .X(_10386_));
 sky130_fd_sc_hd__mux2_1 _15812_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net262),
    .X(_10387_));
 sky130_fd_sc_hd__a221o_1 _15813_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(net3764),
    .B1(_10387_),
    .B2(net3885),
    .C1(net294),
    .X(_10388_));
 sky130_fd_sc_hd__o211ai_1 _15814_ (.A1(net3817),
    .A2(_10386_),
    .B1(_10388_),
    .C1(net3762),
    .Y(_10389_));
 sky130_fd_sc_hd__o311a_4 _15815_ (.A1(net3846),
    .A2(net3812),
    .A3(_10375_),
    .B1(_10385_),
    .C1(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_974 ();
 sky130_fd_sc_hd__o211ai_1 _15817_ (.A1(_08355_),
    .A2(_08735_),
    .B1(net3836),
    .C1(_08348_),
    .Y(_10392_));
 sky130_fd_sc_hd__o21ai_4 _15818_ (.A1(_08348_),
    .A2(_10390_),
    .B1(_10392_),
    .Y(_10393_));
 sky130_fd_sc_hd__mux4_2 _15819_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net3934),
    .S1(net3915),
    .X(_10394_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(net3901),
    .B(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__mux2i_1 _15821_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net3933),
    .Y(_10396_));
 sky130_fd_sc_hd__a21oi_1 _15822_ (.A1(net3933),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .B1(net3914),
    .Y(_10397_));
 sky130_fd_sc_hd__a211o_1 _15823_ (.A1(net3914),
    .A2(_10396_),
    .B1(_10397_),
    .C1(net3901),
    .X(_10398_));
 sky130_fd_sc_hd__mux4_2 _15824_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net267),
    .S1(net3916),
    .X(_10399_));
 sky130_fd_sc_hd__mux4_2 _15825_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net267),
    .S1(net3916),
    .X(_10400_));
 sky130_fd_sc_hd__mux2i_2 _15826_ (.A0(_10399_),
    .A1(_10400_),
    .S(_08109_),
    .Y(_10401_));
 sky130_fd_sc_hd__a32oi_4 _15827_ (.A1(net3781),
    .A2(_10395_),
    .A3(_10398_),
    .B1(_10401_),
    .B2(_08694_),
    .Y(_10402_));
 sky130_fd_sc_hd__mux2i_1 _15828_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .S(net3934),
    .Y(_10403_));
 sky130_fd_sc_hd__mux2i_1 _15829_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .S(net3934),
    .Y(_10404_));
 sky130_fd_sc_hd__a22oi_1 _15830_ (.A1(net3793),
    .A2(_10403_),
    .B1(_10404_),
    .B2(net3775),
    .Y(_10405_));
 sky130_fd_sc_hd__mux2i_1 _15831_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S(net3934),
    .Y(_10406_));
 sky130_fd_sc_hd__mux2i_1 _15832_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S(net3934),
    .Y(_10407_));
 sky130_fd_sc_hd__a22oi_1 _15833_ (.A1(net3780),
    .A2(_10406_),
    .B1(_10407_),
    .B2(net3791),
    .Y(_10408_));
 sky130_fd_sc_hd__a21o_4 _15834_ (.A1(_10405_),
    .A2(_10408_),
    .B1(net3768),
    .X(_10409_));
 sky130_fd_sc_hd__mux4_2 _15835_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S0(net267),
    .S1(net3915),
    .X(_10410_));
 sky130_fd_sc_hd__nand2_2 _15836_ (.A(net3901),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__mux4_2 _15837_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S0(net267),
    .S1(net3915),
    .X(_10412_));
 sky130_fd_sc_hd__nand2_1 _15838_ (.A(_08109_),
    .B(_10412_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand3_4 _15839_ (.A(net3773),
    .B(_10411_),
    .C(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__nand3_4 _15840_ (.A(_10402_),
    .B(_10409_),
    .C(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_973 ();
 sky130_fd_sc_hd__o22ai_1 _15842_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .B2(net3786),
    .Y(_10417_));
 sky130_fd_sc_hd__a221oi_1 _15843_ (.A1(net3736),
    .A2(_10390_),
    .B1(net3675),
    .B2(net3949),
    .C1(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_972 ();
 sky130_fd_sc_hd__o22ai_1 _15845_ (.A1(net3626),
    .A2(_10393_),
    .B1(_10418_),
    .B2(net3747),
    .Y(_10420_));
 sky130_fd_sc_hd__a21oi_1 _15846_ (.A1(net3624),
    .A2(_10393_),
    .B1(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__inv_4 _15847_ (.A(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .Y(_10422_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_971 ();
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(net3722),
    .B(_10415_),
    .Y(_10424_));
 sky130_fd_sc_hd__a21oi_1 _15850_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net3722),
    .B1(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__nand2_2 _15851_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(net3665),
    .Y(_10426_));
 sky130_fd_sc_hd__o21ai_4 _15852_ (.A1(net3666),
    .A2(_10425_),
    .B1(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__nand2_1 _15853_ (.A(net3745),
    .B(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__o31ai_1 _15854_ (.A1(_10422_),
    .A2(net3737),
    .A3(_08171_),
    .B1(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__xnor2_1 _15855_ (.A(_10421_),
    .B(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__mux4_2 _15856_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net3933),
    .S1(net3914),
    .X(_10431_));
 sky130_fd_sc_hd__mux4_2 _15857_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net3918),
    .S1(net3906),
    .X(_10432_));
 sky130_fd_sc_hd__o22ai_1 _15858_ (.A1(net3768),
    .A2(_10431_),
    .B1(_10432_),
    .B2(net3769),
    .Y(_10433_));
 sky130_fd_sc_hd__nand2_1 _15859_ (.A(net3901),
    .B(_10433_),
    .Y(_10434_));
 sky130_fd_sc_hd__mux4_2 _15860_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net3933),
    .S1(net3914),
    .X(_10435_));
 sky130_fd_sc_hd__mux4_2 _15861_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S0(net3918),
    .S1(net3906),
    .X(_10436_));
 sky130_fd_sc_hd__o22ai_1 _15862_ (.A1(net3768),
    .A2(_10435_),
    .B1(_10436_),
    .B2(net3769),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_08109_),
    .B(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__mux2_1 _15864_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net3933),
    .X(_10439_));
 sky130_fd_sc_hd__a22oi_1 _15865_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A2(net3789),
    .B1(_10439_),
    .B2(net3914),
    .Y(_10440_));
 sky130_fd_sc_hd__mux4_2 _15866_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net3933),
    .S1(net3914),
    .X(_10441_));
 sky130_fd_sc_hd__nand2_1 _15867_ (.A(net3901),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__o211ai_1 _15868_ (.A1(net3901),
    .A2(_10440_),
    .B1(_10442_),
    .C1(net3781),
    .Y(_10443_));
 sky130_fd_sc_hd__mux4_2 _15869_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net3918),
    .S1(net3906),
    .X(_10444_));
 sky130_fd_sc_hd__mux4_2 _15870_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net3918),
    .S1(net3906),
    .X(_10445_));
 sky130_fd_sc_hd__mux2i_1 _15871_ (.A0(_10444_),
    .A1(_10445_),
    .S(_08109_),
    .Y(_10446_));
 sky130_fd_sc_hd__nand2_1 _15872_ (.A(_08694_),
    .B(_10446_),
    .Y(_10447_));
 sky130_fd_sc_hd__nand4_1 _15873_ (.A(_10434_),
    .B(_10438_),
    .C(_10443_),
    .D(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(net3722),
    .B(net3674),
    .Y(_10449_));
 sky130_fd_sc_hd__a21oi_2 _15875_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net3722),
    .B1(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__nand2_2 _15876_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(net3665),
    .Y(_10451_));
 sky130_fd_sc_hd__o21a_4 _15877_ (.A1(net3666),
    .A2(_10450_),
    .B1(_10451_),
    .X(_10452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_970 ();
 sky130_fd_sc_hd__a21oi_1 _15879_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(_07864_),
    .B1(net3745),
    .Y(_10454_));
 sky130_fd_sc_hd__a21oi_2 _15880_ (.A1(net3745),
    .A2(_10452_),
    .B1(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__mux4_2 _15881_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net3895),
    .S1(net359),
    .X(_10456_));
 sky130_fd_sc_hd__mux2i_1 _15882_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net3866),
    .Y(_10457_));
 sky130_fd_sc_hd__o2bb2ai_1 _15883_ (.A1_N(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A2_N(net3764),
    .B1(_10457_),
    .B2(_07935_),
    .Y(_10458_));
 sky130_fd_sc_hd__mux4_2 _15884_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net3881),
    .S1(net3862),
    .X(_10459_));
 sky130_fd_sc_hd__mux4_2 _15885_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net3895),
    .S1(net3862),
    .X(_10460_));
 sky130_fd_sc_hd__mux4_2 _15886_ (.A0(_10456_),
    .A1(_10458_),
    .A2(_10459_),
    .A3(_10460_),
    .S0(_07927_),
    .S1(net3848),
    .X(_10461_));
 sky130_fd_sc_hd__mux4_2 _15887_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net3862),
    .S1(net3851),
    .X(_10462_));
 sky130_fd_sc_hd__nand2_2 _15888_ (.A(net3881),
    .B(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__mux4_2 _15889_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .S0(net3862),
    .S1(net3851),
    .X(_10464_));
 sky130_fd_sc_hd__nand2_2 _15890_ (.A(_07935_),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand4_1 _15891_ (.A(net3845),
    .B(net3812),
    .C(_10463_),
    .D(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__mux2i_1 _15892_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S(net3862),
    .Y(_10467_));
 sky130_fd_sc_hd__mux2_1 _15893_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S(net3862),
    .X(_10468_));
 sky130_fd_sc_hd__a21oi_1 _15894_ (.A1(net3803),
    .A2(_10468_),
    .B1(_08839_),
    .Y(_10469_));
 sky130_fd_sc_hd__mux4_2 _15895_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net3862),
    .S1(net3851),
    .X(_10470_));
 sky130_fd_sc_hd__mux4_2 _15896_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .S0(net3862),
    .S1(net3851),
    .X(_10471_));
 sky130_fd_sc_hd__o21ai_0 _15897_ (.A1(_07935_),
    .A2(_10470_),
    .B1(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__o211ai_1 _15898_ (.A1(net3814),
    .A2(_10467_),
    .B1(_10469_),
    .C1(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__o211a_4 _15899_ (.A1(net3845),
    .A2(_10461_),
    .B1(_10466_),
    .C1(_10473_),
    .X(_10474_));
 sky130_fd_sc_hd__o22ai_1 _15900_ (.A1(_08169_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .B2(net3786),
    .Y(_10475_));
 sky130_fd_sc_hd__a21oi_1 _15901_ (.A1(net3949),
    .A2(net3674),
    .B1(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__o21ai_0 _15902_ (.A1(_08172_),
    .A2(_10474_),
    .B1(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__a21oi_1 _15903_ (.A1(net3837),
    .A2(net316),
    .B1(_09680_),
    .Y(_10478_));
 sky130_fd_sc_hd__nand2_2 _15904_ (.A(net3728),
    .B(_10474_),
    .Y(_10479_));
 sky130_fd_sc_hd__o21ai_4 _15905_ (.A1(net3728),
    .A2(_10478_),
    .B1(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__nor2_1 _15906_ (.A(net3626),
    .B(_10480_),
    .Y(_10481_));
 sky130_fd_sc_hd__a221o_4 _15907_ (.A1(net3756),
    .A2(_10477_),
    .B1(_10480_),
    .B2(net3624),
    .C1(_10481_),
    .X(_10482_));
 sky130_fd_sc_hd__nor2_1 _15908_ (.A(_10455_),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__and2_0 _15909_ (.A(_10272_),
    .B(_10302_),
    .X(_10484_));
 sky130_fd_sc_hd__nand2_1 _15910_ (.A(_10338_),
    .B(_10369_),
    .Y(_10485_));
 sky130_fd_sc_hd__o21ai_0 _15911_ (.A1(_10272_),
    .A2(_10302_),
    .B1(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__inv_1 _15912_ (.A(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__nor2_1 _15913_ (.A(_10338_),
    .B(_10369_),
    .Y(_10488_));
 sky130_fd_sc_hd__a221oi_4 _15914_ (.A1(_10484_),
    .A2(_10485_),
    .B1(_10307_),
    .B2(_10487_),
    .C1(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__nand2_1 _15915_ (.A(_10455_),
    .B(_10482_),
    .Y(_10490_));
 sky130_fd_sc_hd__o21ai_1 _15916_ (.A1(_10483_),
    .A2(_10489_),
    .B1(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__xnor2_1 _15917_ (.A(_10430_),
    .B(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__inv_6 _15918_ (.A(net3471),
    .Y(net173));
 sky130_fd_sc_hd__xor2_1 _15919_ (.A(_10455_),
    .B(_10482_),
    .X(_10493_));
 sky130_fd_sc_hd__xnor2_2 _15920_ (.A(net479),
    .B(_10493_),
    .Y(net172));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_969 ();
 sky130_fd_sc_hd__inv_8 _15922_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_10495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_967 ();
 sky130_fd_sc_hd__nor2b_4 _15925_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B_N(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Y(_10498_));
 sky130_fd_sc_hd__and2_4 _15926_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .B(_10498_),
    .X(_10499_));
 sky130_fd_sc_hd__nand2_8 _15927_ (.A(_10495_),
    .B(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__inv_4 _15928_ (.A(\cs_registers_i.debug_mode_i ),
    .Y(_10501_));
 sky130_fd_sc_hd__nor2b_4 _15929_ (.A(net3848),
    .B_N(net366),
    .Y(_10502_));
 sky130_fd_sc_hd__nand4_1 _15930_ (.A(net3858),
    .B(net3839),
    .C(net3804),
    .D(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__nand3_4 _15931_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(net3750),
    .C(net3785),
    .Y(_10504_));
 sky130_fd_sc_hd__or2_4 _15932_ (.A(_10503_),
    .B(_10504_),
    .X(_10505_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(net348),
    .B(net355),
    .Y(_10506_));
 sky130_fd_sc_hd__nor3_4 _15934_ (.A(_07958_),
    .B(_08013_),
    .C(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__nand2_4 _15935_ (.A(net3797),
    .B(_10507_),
    .Y(_10508_));
 sky130_fd_sc_hd__nor2_1 _15936_ (.A(_10505_),
    .B(_10508_),
    .Y(_10509_));
 sky130_fd_sc_hd__nor2_4 _15937_ (.A(net3938),
    .B(net3941),
    .Y(_10510_));
 sky130_fd_sc_hd__nor4_4 _15938_ (.A(net3845),
    .B(net379),
    .C(net3841),
    .D(net354),
    .Y(_10511_));
 sky130_fd_sc_hd__nand2_8 _15939_ (.A(net3797),
    .B(_10511_),
    .Y(_10512_));
 sky130_fd_sc_hd__nand2_1 _15940_ (.A(net3803),
    .B(_10502_),
    .Y(_10513_));
 sky130_fd_sc_hd__or4_4 _15941_ (.A(net3858),
    .B(net3839),
    .C(_10512_),
    .D(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__o21ai_4 _15942_ (.A1(_10507_),
    .A2(_10511_),
    .B1(net3797),
    .Y(_10515_));
 sky130_fd_sc_hd__a21oi_2 _15943_ (.A1(_10503_),
    .A2(_10514_),
    .B1(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__nor4_4 _15944_ (.A(net3858),
    .B(net3851),
    .C(net380),
    .D(_09038_),
    .Y(_10517_));
 sky130_fd_sc_hd__nor4_4 _15945_ (.A(net3901),
    .B(net3915),
    .C(net3933),
    .D(_08538_),
    .Y(_10518_));
 sky130_fd_sc_hd__nor3_4 _15946_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .Y(_10519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_966 ();
 sky130_fd_sc_hd__nor3_1 _15948_ (.A(net3935),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .Y(_10521_));
 sky130_fd_sc_hd__o2111ai_2 _15949_ (.A1(_10516_),
    .A2(_10517_),
    .B1(_10518_),
    .C1(_10519_),
    .D1(_10521_),
    .Y(_10522_));
 sky130_fd_sc_hd__a21oi_1 _15950_ (.A1(net3939),
    .A2(_08019_),
    .B1(_08014_),
    .Y(_10523_));
 sky130_fd_sc_hd__o221ai_2 _15951_ (.A1(net3842),
    .A2(_08021_),
    .B1(net381),
    .B2(_10523_),
    .C1(_08028_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand3_2 _15952_ (.A(_08033_),
    .B(_08073_),
    .C(_08006_),
    .Y(_10525_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(net3830),
    .B(_07906_),
    .Y(_10526_));
 sky130_fd_sc_hd__o21ai_0 _15954_ (.A1(_08081_),
    .A2(_08003_),
    .B1(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__a311oi_1 _15955_ (.A1(net3938),
    .A2(_07883_),
    .A3(_10527_),
    .B1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .C1(_08048_),
    .Y(_10528_));
 sky130_fd_sc_hd__a21oi_1 _15956_ (.A1(net3938),
    .A2(net3941),
    .B1(net3935),
    .Y(_10529_));
 sky130_fd_sc_hd__nor2_1 _15957_ (.A(_08038_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__nor2_1 _15958_ (.A(net3838),
    .B(_08184_),
    .Y(_10531_));
 sky130_fd_sc_hd__o21bai_1 _15959_ (.A1(_07879_),
    .A2(_10531_),
    .B1_N(net3835),
    .Y(_10532_));
 sky130_fd_sc_hd__o32ai_1 _15960_ (.A1(net330),
    .A2(_07884_),
    .A3(net3785),
    .B1(_08025_),
    .B2(_07897_),
    .Y(_10533_));
 sky130_fd_sc_hd__a222oi_1 _15961_ (.A1(net3753),
    .A2(_10530_),
    .B1(_10532_),
    .B2(_08186_),
    .C1(_10533_),
    .C2(_07895_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand4_1 _15962_ (.A(_10524_),
    .B(_10525_),
    .C(_10528_),
    .D(_10534_),
    .Y(_10535_));
 sky130_fd_sc_hd__a31oi_4 _15963_ (.A1(_08188_),
    .A2(_10510_),
    .A3(_10522_),
    .B1(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_965 ();
 sky130_fd_sc_hd__nand2b_4 _15965_ (.A_N(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_10538_));
 sky130_fd_sc_hd__nor2_4 _15966_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__nand2_8 _15967_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10539_),
    .Y(_10540_));
 sky130_fd_sc_hd__nor3b_4 _15968_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(_10540_),
    .C_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_10541_));
 sky130_fd_sc_hd__and2_4 _15969_ (.A(net3612),
    .B(_10541_),
    .X(_10542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_963 ();
 sky130_fd_sc_hd__a211oi_4 _15972_ (.A1(net356),
    .A2(_10518_),
    .B1(_10510_),
    .C1(_08405_),
    .Y(_10545_));
 sky130_fd_sc_hd__nand2_8 _15973_ (.A(_10542_),
    .B(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__mux2i_4 _15974_ (.A0(net3707),
    .A1(_08736_),
    .S(net3718),
    .Y(_10547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_962 ();
 sky130_fd_sc_hd__nand2_8 _15976_ (.A(net3738),
    .B(_10536_),
    .Y(_10549_));
 sky130_fd_sc_hd__a41oi_4 _15977_ (.A1(net3749),
    .A2(_08348_),
    .A3(_08447_),
    .A4(_08448_),
    .B1(_08489_),
    .Y(_10550_));
 sky130_fd_sc_hd__nor2_4 _15978_ (.A(_08359_),
    .B(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__nor2_2 _15979_ (.A(_10549_),
    .B(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__nand2_2 _15980_ (.A(net3586),
    .B(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__nand2b_4 _15981_ (.A_N(_08000_),
    .B(_08779_),
    .Y(_10554_));
 sky130_fd_sc_hd__and3_4 _15982_ (.A(_08241_),
    .B(net3738),
    .C(_10536_),
    .X(_10555_));
 sky130_fd_sc_hd__nand2b_4 _15983_ (.A_N(_10554_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__and2_4 _15984_ (.A(_08406_),
    .B(_10536_),
    .X(_10557_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_961 ();
 sky130_fd_sc_hd__nand4_1 _15986_ (.A(net3618),
    .B(_08919_),
    .C(net3614),
    .D(_10557_),
    .Y(_10559_));
 sky130_fd_sc_hd__nor2_4 _15987_ (.A(net353),
    .B(_10549_),
    .Y(_10560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_960 ();
 sky130_fd_sc_hd__nand2_1 _15989_ (.A(_08737_),
    .B(_10557_),
    .Y(_10562_));
 sky130_fd_sc_hd__inv_4 _15990_ (.A(net3614),
    .Y(_10563_));
 sky130_fd_sc_hd__nand4_1 _15991_ (.A(net3618),
    .B(net3616),
    .C(_10563_),
    .D(_10557_),
    .Y(_10564_));
 sky130_fd_sc_hd__or4_4 _15992_ (.A(_10556_),
    .B(_10560_),
    .C(_10562_),
    .D(_10564_),
    .X(_10565_));
 sky130_fd_sc_hd__nand2_8 _15993_ (.A(net3623),
    .B(net3622),
    .Y(_10566_));
 sky130_fd_sc_hd__nand2_8 _15994_ (.A(_10557_),
    .B(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__nand2b_4 _15995_ (.A_N(_10565_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__o31ai_1 _15996_ (.A1(_09026_),
    .A2(_10556_),
    .A3(_10559_),
    .B1(_10568_),
    .Y(_10569_));
 sky130_fd_sc_hd__or2_4 _15997_ (.A(_08000_),
    .B(_08779_),
    .X(_10570_));
 sky130_fd_sc_hd__nand2_4 _15998_ (.A(_09026_),
    .B(_10557_),
    .Y(_10571_));
 sky130_fd_sc_hd__nor2_4 _15999_ (.A(_10570_),
    .B(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_958 ();
 sky130_fd_sc_hd__nor3_4 _16002_ (.A(net3621),
    .B(net308),
    .C(_10549_),
    .Y(_10575_));
 sky130_fd_sc_hd__nand2_8 _16003_ (.A(_10551_),
    .B(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__nor2_4 _16004_ (.A(_08737_),
    .B(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__nor3_4 _16005_ (.A(_08241_),
    .B(_10577_),
    .C(_10559_),
    .Y(_10578_));
 sky130_fd_sc_hd__and2_4 _16006_ (.A(_10572_),
    .B(_10578_),
    .X(_10579_));
 sky130_fd_sc_hd__nor2_4 _16007_ (.A(_10554_),
    .B(_10571_),
    .Y(_10580_));
 sky130_fd_sc_hd__and2_4 _16008_ (.A(_10580_),
    .B(_10578_),
    .X(_10581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_957 ();
 sky130_fd_sc_hd__nor2_4 _16010_ (.A(_10579_),
    .B(_10581_),
    .Y(_10583_));
 sky130_fd_sc_hd__o21ai_4 _16011_ (.A1(net3619),
    .A2(net3595),
    .B1(_10557_),
    .Y(_10584_));
 sky130_fd_sc_hd__nand2_8 _16012_ (.A(_10567_),
    .B(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__nor2_4 _16013_ (.A(_08241_),
    .B(_08737_),
    .Y(_10586_));
 sky130_fd_sc_hd__nand2_4 _16014_ (.A(_08000_),
    .B(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nor2_2 _16015_ (.A(_08779_),
    .B(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__nor2_4 _16016_ (.A(_09026_),
    .B(_10559_),
    .Y(_10589_));
 sky130_fd_sc_hd__nand2_8 _16017_ (.A(_10588_),
    .B(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__nor2_2 _16018_ (.A(_10585_),
    .B(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__nor2_1 _16019_ (.A(_08000_),
    .B(_08779_),
    .Y(_10592_));
 sky130_fd_sc_hd__a21oi_2 _16020_ (.A1(_10592_),
    .A2(_10586_),
    .B1(_10549_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand2b_4 _16021_ (.A_N(_10593_),
    .B(_10589_),
    .Y(_10594_));
 sky130_fd_sc_hd__nor2_4 _16022_ (.A(_10585_),
    .B(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__nand2_4 _16023_ (.A(_10547_),
    .B(_10551_),
    .Y(_10596_));
 sky130_fd_sc_hd__a21oi_2 _16024_ (.A1(net3619),
    .A2(net3595),
    .B1(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_1 _16025_ (.A(_10555_),
    .B(_10589_),
    .Y(_10598_));
 sky130_fd_sc_hd__nor3_1 _16026_ (.A(_10570_),
    .B(_10597_),
    .C(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__nor2_4 _16027_ (.A(net3619),
    .B(net308),
    .Y(_10600_));
 sky130_fd_sc_hd__nor2_4 _16028_ (.A(_08359_),
    .B(_08490_),
    .Y(_10601_));
 sky130_fd_sc_hd__nand3_4 _16029_ (.A(_10557_),
    .B(_10600_),
    .C(_10601_),
    .Y(_10602_));
 sky130_fd_sc_hd__nand2b_4 _16030_ (.A_N(_10602_),
    .B(_10572_),
    .Y(_10603_));
 sky130_fd_sc_hd__nor4_2 _16031_ (.A(_08241_),
    .B(_10603_),
    .C(_10562_),
    .D(_10564_),
    .Y(_10604_));
 sky130_fd_sc_hd__nor4_1 _16032_ (.A(_10591_),
    .B(_10595_),
    .C(_10599_),
    .D(_10604_),
    .Y(_10605_));
 sky130_fd_sc_hd__nor2_1 _16033_ (.A(_10576_),
    .B(_10594_),
    .Y(_10606_));
 sky130_fd_sc_hd__a2111oi_1 _16034_ (.A1(_10557_),
    .A2(_10570_),
    .B1(_10585_),
    .C1(_10598_),
    .D1(_08737_),
    .Y(_10607_));
 sky130_fd_sc_hd__nor2_1 _16035_ (.A(_10606_),
    .B(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__nand3_1 _16036_ (.A(_10583_),
    .B(_10605_),
    .C(_10608_),
    .Y(_10609_));
 sky130_fd_sc_hd__and3_4 _16037_ (.A(net3621),
    .B(net3595),
    .C(_10557_),
    .X(_10610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_956 ();
 sky130_fd_sc_hd__nand2_4 _16039_ (.A(_10567_),
    .B(_10610_),
    .Y(_10612_));
 sky130_fd_sc_hd__nor2_4 _16040_ (.A(_10612_),
    .B(_10590_),
    .Y(_10613_));
 sky130_fd_sc_hd__nand2_2 _16041_ (.A(_10575_),
    .B(_10601_),
    .Y(_10614_));
 sky130_fd_sc_hd__nor2_2 _16042_ (.A(_10614_),
    .B(_10594_),
    .Y(_10615_));
 sky130_fd_sc_hd__and2_4 _16043_ (.A(net308),
    .B(_10557_),
    .X(_10616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_955 ();
 sky130_fd_sc_hd__nand3_2 _16045_ (.A(net3619),
    .B(_10551_),
    .C(_10616_),
    .Y(_10618_));
 sky130_fd_sc_hd__nor2_2 _16046_ (.A(_10618_),
    .B(_10590_),
    .Y(_10619_));
 sky130_fd_sc_hd__nor2_4 _16047_ (.A(_10602_),
    .B(_10594_),
    .Y(_10620_));
 sky130_fd_sc_hd__or4_4 _16048_ (.A(_10613_),
    .B(_10615_),
    .C(_10619_),
    .D(_10620_),
    .X(_10621_));
 sky130_fd_sc_hd__nor2_2 _16049_ (.A(_10552_),
    .B(_10560_),
    .Y(_10622_));
 sky130_fd_sc_hd__nor3_1 _16050_ (.A(_10587_),
    .B(_10616_),
    .C(_10564_),
    .Y(_10623_));
 sky130_fd_sc_hd__nor2_4 _16051_ (.A(_10602_),
    .B(_10590_),
    .Y(_10624_));
 sky130_fd_sc_hd__nor2_4 _16052_ (.A(_10576_),
    .B(_10590_),
    .Y(_10625_));
 sky130_fd_sc_hd__a311o_1 _16053_ (.A1(_08779_),
    .A2(_10622_),
    .A3(_10623_),
    .B1(_10624_),
    .C1(_10625_),
    .X(_10626_));
 sky130_fd_sc_hd__a2111oi_2 _16054_ (.A1(_10553_),
    .A2(_10569_),
    .B1(_10609_),
    .C1(_10621_),
    .D1(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_953 ();
 sky130_fd_sc_hd__inv_1 _16057_ (.A(\cs_registers_i.priv_mode_id_o[0] ),
    .Y(_10630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_952 ();
 sky130_fd_sc_hd__a21oi_1 _16059_ (.A1(_10630_),
    .A2(net3616),
    .B1(net3618),
    .Y(_10632_));
 sky130_fd_sc_hd__nor2_1 _16060_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__a31oi_1 _16061_ (.A1(_10630_),
    .A2(net3618),
    .A3(net3616),
    .B1(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__or2_4 _16062_ (.A(_10549_),
    .B(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__o21ai_2 _16063_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10568_),
    .B1(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__nor2_2 _16064_ (.A(_10627_),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__o31ai_4 _16065_ (.A1(net353),
    .A2(net3614),
    .A3(_10546_),
    .B1(_10637_),
    .Y(_10638_));
 sky130_fd_sc_hd__nand2_8 _16066_ (.A(net3738),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__nand2_2 _16067_ (.A(net3612),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__nor2_1 _16068_ (.A(_10504_),
    .B(_10514_),
    .Y(_10641_));
 sky130_fd_sc_hd__nor2_4 _16069_ (.A(_10505_),
    .B(_10512_),
    .Y(_10642_));
 sky130_fd_sc_hd__a21oi_1 _16070_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_10641_),
    .B1(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__a21oi_1 _16071_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(net3950),
    .B1(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__a221o_1 _16072_ (.A1(_10501_),
    .A2(_10509_),
    .B1(_10640_),
    .B2(\id_stage_i.controller_i.instr_valid_i ),
    .C1(_10644_),
    .X(_10645_));
 sky130_fd_sc_hd__and2_0 _16073_ (.A(_10500_),
    .B(_10645_),
    .X(\id_stage_i.controller_i.illegal_insn_d ));
 sky130_fd_sc_hd__nand2_8 _16074_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Y(_10646_));
 sky130_fd_sc_hd__nand2b_4 _16075_ (.A_N(_10504_),
    .B(_10517_),
    .Y(_10647_));
 sky130_fd_sc_hd__nand2_2 _16076_ (.A(_10646_),
    .B(_10647_),
    .Y(_10648_));
 sky130_fd_sc_hd__or2_4 _16077_ (.A(_10645_),
    .B(_10648_),
    .X(_10649_));
 sky130_fd_sc_hd__nand2_2 _16078_ (.A(_10500_),
    .B(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__inv_1 _16079_ (.A(_10650_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 sky130_fd_sc_hd__inv_1 _16080_ (.A(\load_store_unit_i.data_we_q ),
    .Y(_10651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_951 ();
 sky130_fd_sc_hd__nor3_4 _16082_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(\load_store_unit_i.ls_fsm_cs[0] ),
    .C(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_10653_));
 sky130_fd_sc_hd__and2_4 _16083_ (.A(net59),
    .B(_10653_),
    .X(_10654_));
 sky130_fd_sc_hd__o21ai_4 _16084_ (.A1(net25),
    .A2(\load_store_unit_i.lsu_err_q ),
    .B1(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__nor2_1 _16085_ (.A(_10651_),
    .B(_10655_),
    .Y(\id_stage_i.controller_i.store_err_i ));
 sky130_fd_sc_hd__nor2_1 _16086_ (.A(\load_store_unit_i.data_we_q ),
    .B(_10655_),
    .Y(\id_stage_i.controller_i.load_err_i ));
 sky130_fd_sc_hd__inv_4 _16087_ (.A(\load_store_unit_i.data_type_q[2] ),
    .Y(_10656_));
 sky130_fd_sc_hd__and2_4 _16088_ (.A(net3753),
    .B(_10536_),
    .X(_10657_));
 sky130_fd_sc_hd__nor2b_4 _16089_ (.A(\id_stage_i.id_fsm_q ),
    .B_N(_10541_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand3_4 _16090_ (.A(_10653_),
    .B(_10657_),
    .C(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__clkinv_2 _16091_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .Y(_10660_));
 sky130_fd_sc_hd__nand2_2 _16092_ (.A(_10660_),
    .B(\load_store_unit_i.ls_fsm_cs[0] ),
    .Y(_10661_));
 sky130_fd_sc_hd__a21boi_4 _16093_ (.A1(_10659_),
    .A2(_10661_),
    .B1_N(net26),
    .Y(_10662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_950 ();
 sky130_fd_sc_hd__nand3_1 _16095_ (.A(net3753),
    .B(_08033_),
    .C(_10662_),
    .Y(_10664_));
 sky130_fd_sc_hd__o21ai_0 _16096_ (.A1(_10656_),
    .A2(_10662_),
    .B1(_10664_),
    .Y(_00007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_949 ();
 sky130_fd_sc_hd__inv_6 _16098_ (.A(\load_store_unit_i.data_type_q[1] ),
    .Y(_10666_));
 sky130_fd_sc_hd__nand3_1 _16099_ (.A(net3753),
    .B(_10510_),
    .C(_10662_),
    .Y(_10667_));
 sky130_fd_sc_hd__o21ai_0 _16100_ (.A1(_10666_),
    .A2(_10662_),
    .B1(_10667_),
    .Y(_00006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_945 ();
 sky130_fd_sc_hd__inv_6 _16105_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_10672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_944 ();
 sky130_fd_sc_hd__nand2_8 _16107_ (.A(_10672_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10674_));
 sky130_fd_sc_hd__nor3_4 _16108_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_10674_),
    .Y(_10675_));
 sky130_fd_sc_hd__nand2b_4 _16109_ (.A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_942 ();
 sky130_fd_sc_hd__nand3_4 _16112_ (.A(net3937),
    .B(net3739),
    .C(_10542_),
    .Y(_10679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_941 ();
 sky130_fd_sc_hd__o21ai_0 _16114_ (.A1(_10676_),
    .A2(_10679_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Y(_10681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_940 ();
 sky130_fd_sc_hd__and3_4 _16116_ (.A(net3937),
    .B(net3739),
    .C(_10542_),
    .X(_10683_));
 sky130_fd_sc_hd__nand2_8 _16117_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_939 ();
 sky130_fd_sc_hd__nand2_1 _16119_ (.A(_10681_),
    .B(_10684_),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_1 _16120_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .Y(_10686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_936 ();
 sky130_fd_sc_hd__nor2_4 _16124_ (.A(_08009_),
    .B(net3747),
    .Y(_10690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_934 ();
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(_10542_),
    .B(net3734),
    .Y(_10693_));
 sky130_fd_sc_hd__nor3_1 _16128_ (.A(net152),
    .B(net151),
    .C(net3514),
    .Y(_10694_));
 sky130_fd_sc_hd__xnor2_1 _16129_ (.A(_08320_),
    .B(net3553),
    .Y(net176));
 sky130_fd_sc_hd__nor2_1 _16130_ (.A(_08413_),
    .B(_08672_),
    .Y(_10695_));
 sky130_fd_sc_hd__xnor2_1 _16131_ (.A(_08711_),
    .B(_08742_),
    .Y(_10696_));
 sky130_fd_sc_hd__xnor2_1 _16132_ (.A(_10695_),
    .B(_10696_),
    .Y(net175));
 sky130_fd_sc_hd__o21ai_0 _16133_ (.A1(net299),
    .A2(net3619),
    .B1(_08627_),
    .Y(_10697_));
 sky130_fd_sc_hd__xor2_1 _16134_ (.A(_08622_),
    .B(_10697_),
    .X(_10698_));
 sky130_fd_sc_hd__xnor2_1 _16135_ (.A(net3621),
    .B(net3620),
    .Y(_10699_));
 sky130_fd_sc_hd__nand2_2 _16136_ (.A(net3744),
    .B(_10699_),
    .Y(_10700_));
 sky130_fd_sc_hd__o21ai_4 _16137_ (.A1(_08498_),
    .A2(_10698_),
    .B1(_10700_),
    .Y(_10701_));
 sky130_fd_sc_hd__o21a_1 _16138_ (.A1(_08497_),
    .A2(net3576),
    .B1(_08671_),
    .X(_10702_));
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B(_07864_),
    .Y(_10703_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(_08401_),
    .B(_08399_),
    .Y(_10704_));
 sky130_fd_sc_hd__xor2_1 _16141_ (.A(_10703_),
    .B(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__xnor2_1 _16142_ (.A(_08205_),
    .B(net3599),
    .Y(_10706_));
 sky130_fd_sc_hd__xnor2_1 _16143_ (.A(net3623),
    .B(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__nor2_1 _16144_ (.A(_07857_),
    .B(_10707_),
    .Y(_10708_));
 sky130_fd_sc_hd__a21oi_1 _16145_ (.A1(_07857_),
    .A2(_10705_),
    .B1(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__xor2_1 _16146_ (.A(_10702_),
    .B(_10709_),
    .X(_10710_));
 sky130_fd_sc_hd__nand2_1 _16147_ (.A(net3626),
    .B(_08490_),
    .Y(_10711_));
 sky130_fd_sc_hd__nand2_1 _16148_ (.A(_08205_),
    .B(_10550_),
    .Y(_10712_));
 sky130_fd_sc_hd__a21oi_1 _16149_ (.A1(_10711_),
    .A2(_10712_),
    .B1(_08494_),
    .Y(_10713_));
 sky130_fd_sc_hd__xnor2_1 _16150_ (.A(net3598),
    .B(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B(_07864_),
    .Y(_10715_));
 sky130_fd_sc_hd__xor2_1 _16152_ (.A(_10715_),
    .B(_08495_),
    .X(_10716_));
 sky130_fd_sc_hd__nand2_2 _16153_ (.A(_07857_),
    .B(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__o21ai_4 _16154_ (.A1(_07857_),
    .A2(_10714_),
    .B1(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__xor2_1 _16155_ (.A(_08547_),
    .B(net3584),
    .X(_10719_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_10718_),
    .B(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__and2_0 _16157_ (.A(_08547_),
    .B(net3584),
    .X(_10721_));
 sky130_fd_sc_hd__nor2_1 _16158_ (.A(_08547_),
    .B(net3584),
    .Y(_10722_));
 sky130_fd_sc_hd__mux2i_1 _16159_ (.A0(_10721_),
    .A1(_10722_),
    .S(_10718_),
    .Y(_10723_));
 sky130_fd_sc_hd__mux2i_1 _16160_ (.A0(_10720_),
    .A1(_10723_),
    .S(net3583),
    .Y(_10724_));
 sky130_fd_sc_hd__nand3_1 _16161_ (.A(_10701_),
    .B(_10710_),
    .C(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__nor4_1 _16162_ (.A(net178),
    .B(net3537),
    .C(net3535),
    .D(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand2_1 _16163_ (.A(_08815_),
    .B(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__or4_4 _16164_ (.A(net180),
    .B(net179),
    .C(net155),
    .D(_10727_),
    .X(_10728_));
 sky130_fd_sc_hd__nor3_1 _16165_ (.A(net156),
    .B(net158),
    .C(_10728_),
    .Y(_10729_));
 sky130_fd_sc_hd__nand3_1 _16166_ (.A(_09945_),
    .B(_10694_),
    .C(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__nor3_1 _16167_ (.A(net157),
    .B(net160),
    .C(net163),
    .Y(_10731_));
 sky130_fd_sc_hd__nand4_1 _16168_ (.A(_09252_),
    .B(_09675_),
    .C(_09812_),
    .D(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__nor4_1 _16169_ (.A(net452),
    .B(net166),
    .C(_10730_),
    .D(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__nor4b_1 _16170_ (.A(net167),
    .B(net170),
    .C(net172),
    .D_N(_10733_),
    .Y(_10734_));
 sky130_fd_sc_hd__nor3_1 _16171_ (.A(net273),
    .B(net168),
    .C(net169),
    .Y(_10735_));
 sky130_fd_sc_hd__and3_4 _16172_ (.A(net3470),
    .B(_10734_),
    .C(_10735_),
    .X(_10736_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(_10679_),
    .Y(_10737_));
 sky130_fd_sc_hd__o31ai_1 _16174_ (.A1(_10686_),
    .A2(_10693_),
    .A3(_10736_),
    .B1(_10737_),
    .Y(_00004_));
 sky130_fd_sc_hd__nand3_4 _16175_ (.A(_08009_),
    .B(net3739),
    .C(_10542_),
    .Y(_10738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_933 ();
 sky130_fd_sc_hd__nand2_8 _16177_ (.A(_08075_),
    .B(_07857_),
    .Y(_10740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_931 ();
 sky130_fd_sc_hd__a21oi_1 _16180_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(_10740_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_1 _16181_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(_10738_),
    .Y(_10744_));
 sky130_fd_sc_hd__o21ai_0 _16182_ (.A1(_10738_),
    .A2(_10743_),
    .B1(_10744_),
    .Y(_00000_));
 sky130_fd_sc_hd__and3_4 _16183_ (.A(_08075_),
    .B(net3820),
    .C(net3819),
    .X(_10745_));
 sky130_fd_sc_hd__and3_4 _16184_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(_08028_),
    .C(_10745_),
    .X(_10746_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_928 ();
 sky130_fd_sc_hd__mux2_1 _16188_ (.A0(_10746_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .S(_10738_),
    .X(_00001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_925 ();
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_10679_),
    .Y(_10753_));
 sky130_fd_sc_hd__o31ai_1 _16193_ (.A1(_07862_),
    .A2(_10676_),
    .A3(_10679_),
    .B1(_10753_),
    .Y(_00002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_923 ();
 sky130_fd_sc_hd__a21oi_1 _16196_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_10736_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_1 _16197_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(_10679_),
    .Y(_10757_));
 sky130_fd_sc_hd__o21ai_0 _16198_ (.A1(_10693_),
    .A2(_10756_),
    .B1(_10757_),
    .Y(_00003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_917 ();
 sky130_fd_sc_hd__mux2i_1 _16205_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10764_));
 sky130_fd_sc_hd__mux2_4 _16206_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10765_));
 sky130_fd_sc_hd__nand2_1 _16207_ (.A(net3948),
    .B(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__o21a_4 _16208_ (.A1(net3948),
    .A2(_10764_),
    .B1(_10766_),
    .X(_10767_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_916 ();
 sky130_fd_sc_hd__inv_16 _16210_ (.A(_10767_),
    .Y(_10769_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_913 ();
 sky130_fd_sc_hd__mux2i_1 _16214_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10772_));
 sky130_fd_sc_hd__mux2_8 _16215_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10773_));
 sky130_fd_sc_hd__nand2_1 _16216_ (.A(net3948),
    .B(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__o21a_4 _16217_ (.A1(net3948),
    .A2(_10772_),
    .B1(_10774_),
    .X(_10775_));
 sky130_fd_sc_hd__inv_16 _16218_ (.A(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_912 ();
 sky130_fd_sc_hd__xnor2_4 _16220_ (.A(net3576),
    .B(_10718_),
    .Y(net171));
 sky130_fd_sc_hd__inv_8 _16221_ (.A(net3533),
    .Y(net174));
 sky130_fd_sc_hd__nor3_2 _16222_ (.A(_10495_),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C(_10538_),
    .Y(_10777_));
 sky130_fd_sc_hd__nor2_1 _16223_ (.A(_07897_),
    .B(_07900_),
    .Y(_10778_));
 sky130_fd_sc_hd__o21ai_2 _16224_ (.A1(_08040_),
    .A2(_10778_),
    .B1(_07895_),
    .Y(_10779_));
 sky130_fd_sc_hd__nand2_4 _16225_ (.A(_10536_),
    .B(_10658_),
    .Y(_10780_));
 sky130_fd_sc_hd__o21bai_4 _16226_ (.A1(_10779_),
    .A2(_10780_),
    .B1_N(\id_stage_i.branch_set ),
    .Y(_10781_));
 sky130_fd_sc_hd__nand2_4 _16227_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .B(_10498_),
    .Y(_10782_));
 sky130_fd_sc_hd__nor2_2 _16228_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10782_),
    .Y(_10783_));
 sky130_fd_sc_hd__or3_4 _16229_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.exc_req_q ),
    .C(\id_stage_i.controller_i.load_err_q ),
    .X(_10784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_910 ();
 sky130_fd_sc_hd__or2_0 _16232_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10647_),
    .X(_10787_));
 sky130_fd_sc_hd__nor2_1 _16233_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(\cs_registers_i.priv_mode_id_o[0] ),
    .Y(_10788_));
 sky130_fd_sc_hd__nand2_1 _16234_ (.A(\cs_registers_i.dcsr_q[12] ),
    .B(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__nand3_1 _16235_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(\cs_registers_i.priv_mode_id_o[0] ),
    .C(\cs_registers_i.dcsr_q[15] ),
    .Y(_10790_));
 sky130_fd_sc_hd__nand2_4 _16236_ (.A(_10789_),
    .B(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__o21ai_0 _16237_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10791_),
    .B1(net3895),
    .Y(_10792_));
 sky130_fd_sc_hd__nor3_1 _16238_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(_10787_),
    .C(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__nand2_2 _16239_ (.A(_10784_),
    .B(_10793_),
    .Y(_10794_));
 sky130_fd_sc_hd__nand2_2 _16240_ (.A(_10783_),
    .B(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__nor2_4 _16241_ (.A(_10505_),
    .B(_10515_),
    .Y(_10796_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_10784_),
    .B(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__nor2_4 _16243_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_10798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_909 ();
 sky130_fd_sc_hd__nor2_1 _16245_ (.A(\cs_registers_i.dcsr_q[2] ),
    .B(net60),
    .Y(_10800_));
 sky130_fd_sc_hd__nand2_1 _16246_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__a21oi_1 _16247_ (.A1(_10798_),
    .A2(_10801_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_10802_));
 sky130_fd_sc_hd__a21oi_2 _16248_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(net147),
    .B1(net145),
    .Y(_10803_));
 sky130_fd_sc_hd__a22o_4 _16249_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net139),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net140),
    .X(_10804_));
 sky130_fd_sc_hd__a22oi_2 _16250_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net141),
    .B1(\cs_registers_i.mie_q[7] ),
    .B2(net142),
    .Y(_10805_));
 sky130_fd_sc_hd__nor2b_4 _16251_ (.A(_10804_),
    .B_N(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__a22oi_2 _16252_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net137),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net138),
    .Y(_10807_));
 sky130_fd_sc_hd__a22oi_2 _16253_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net130),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net136),
    .Y(_10808_));
 sky130_fd_sc_hd__nand3_4 _16254_ (.A(_10806_),
    .B(_10807_),
    .C(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_2 _16255_ (.A(\cs_registers_i.mie_q[12] ),
    .B(net133),
    .Y(_10810_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(\cs_registers_i.mie_q[13] ),
    .B(net134),
    .Y(_10811_));
 sky130_fd_sc_hd__a22oi_2 _16257_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net131),
    .B1(\cs_registers_i.mie_q[11] ),
    .B2(net132),
    .Y(_10812_));
 sky130_fd_sc_hd__and2_4 _16258_ (.A(\cs_registers_i.mie_q[8] ),
    .B(net143),
    .X(_10813_));
 sky130_fd_sc_hd__a21oi_4 _16259_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(net144),
    .B1(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand4_1 _16260_ (.A(_10810_),
    .B(_10811_),
    .C(_10812_),
    .D(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand2_8 _16261_ (.A(\cs_registers_i.mie_q[14] ),
    .B(net135),
    .Y(_10816_));
 sky130_fd_sc_hd__nor3b_4 _16262_ (.A(_10809_),
    .B(_10815_),
    .C_N(_10816_),
    .Y(_10817_));
 sky130_fd_sc_hd__nand2_1 _16263_ (.A(net129),
    .B(\cs_registers_i.mie_q[15] ),
    .Y(_10818_));
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(\cs_registers_i.mie_q[17] ),
    .B(net146),
    .Y(_10819_));
 sky130_fd_sc_hd__and3_4 _16265_ (.A(_10817_),
    .B(_10818_),
    .C(_10819_),
    .X(_10820_));
 sky130_fd_sc_hd__nand2_8 _16266_ (.A(_10803_),
    .B(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__inv_4 _16267_ (.A(\cs_registers_i.nmi_mode_i ),
    .Y(_10822_));
 sky130_fd_sc_hd__o2111a_4 _16268_ (.A1(net145),
    .A2(\cs_registers_i.csr_mstatus_mie_o ),
    .B1(_10821_),
    .C1(_10822_),
    .D1(_10501_),
    .X(_10823_));
 sky130_fd_sc_hd__a21oi_1 _16269_ (.A1(_10499_),
    .A2(_10823_),
    .B1(_10798_),
    .Y(_10824_));
 sky130_fd_sc_hd__o22ai_2 _16270_ (.A1(_10795_),
    .A2(_10797_),
    .B1(_10802_),
    .B2(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__a31o_4 _16271_ (.A1(_10777_),
    .A2(_10646_),
    .A3(_10781_),
    .B1(_10825_),
    .X(_10826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_903 ();
 sky130_fd_sc_hd__o21a_4 _16278_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .A2(net3567),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 sky130_fd_sc_hd__mux2_8 _16279_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_901 ();
 sky130_fd_sc_hd__mux2i_1 _16282_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10836_));
 sky130_fd_sc_hd__nor2_1 _16283_ (.A(net3948),
    .B(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__a21oi_4 _16284_ (.A1(net3948),
    .A2(_10833_),
    .B1(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__inv_2 _16285_ (.A(_10838_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[6] ));
 sky130_fd_sc_hd__mux2i_1 _16286_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10839_));
 sky130_fd_sc_hd__mux2_4 _16287_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10840_));
 sky130_fd_sc_hd__nand2_1 _16288_ (.A(net3948),
    .B(_10840_),
    .Y(_10841_));
 sky130_fd_sc_hd__o21a_4 _16289_ (.A1(net3948),
    .A2(_10839_),
    .B1(_10841_),
    .X(_10842_));
 sky130_fd_sc_hd__inv_6 _16290_ (.A(_10842_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[5] ));
 sky130_fd_sc_hd__mux2i_1 _16291_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10843_));
 sky130_fd_sc_hd__mux2_1 _16292_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10844_));
 sky130_fd_sc_hd__nand2_1 _16293_ (.A(net3948),
    .B(_10844_),
    .Y(_10845_));
 sky130_fd_sc_hd__o21a_4 _16294_ (.A1(net3948),
    .A2(_10843_),
    .B1(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__clkinv_2 _16295_ (.A(_10846_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[7] ));
 sky130_fd_sc_hd__mux2i_1 _16296_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10847_));
 sky130_fd_sc_hd__mux2_4 _16297_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10848_));
 sky130_fd_sc_hd__nand2_1 _16298_ (.A(net3948),
    .B(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__o21ai_4 _16299_ (.A1(net3948),
    .A2(_10847_),
    .B1(_10849_),
    .Y(_10850_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_900 ();
 sky130_fd_sc_hd__mux2i_1 _16301_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10851_));
 sky130_fd_sc_hd__mux2_1 _16302_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10852_));
 sky130_fd_sc_hd__nand2_1 _16303_ (.A(net3948),
    .B(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__o21a_4 _16304_ (.A1(net3948),
    .A2(_10851_),
    .B1(_10853_),
    .X(_10854_));
 sky130_fd_sc_hd__inv_4 _16305_ (.A(_10854_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[9] ));
 sky130_fd_sc_hd__mux2i_1 _16306_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10855_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10856_));
 sky130_fd_sc_hd__nand2_1 _16308_ (.A(net3948),
    .B(_10856_),
    .Y(_10857_));
 sky130_fd_sc_hd__o21a_4 _16309_ (.A1(net3948),
    .A2(_10855_),
    .B1(_10857_),
    .X(_10858_));
 sky130_fd_sc_hd__inv_6 _16310_ (.A(_10858_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[10] ));
 sky130_fd_sc_hd__mux2i_1 _16311_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10859_));
 sky130_fd_sc_hd__mux2_4 _16312_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10860_));
 sky130_fd_sc_hd__nand2_1 _16313_ (.A(net3948),
    .B(_10860_),
    .Y(_10861_));
 sky130_fd_sc_hd__o21ai_4 _16314_ (.A1(net3948),
    .A2(_10859_),
    .B1(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_899 ();
 sky130_fd_sc_hd__mux2i_1 _16316_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10863_));
 sky130_fd_sc_hd__mux2_1 _16317_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10864_));
 sky130_fd_sc_hd__nand2_1 _16318_ (.A(net3948),
    .B(_10864_),
    .Y(_10865_));
 sky130_fd_sc_hd__o21a_4 _16319_ (.A1(net3948),
    .A2(_10863_),
    .B1(_10865_),
    .X(_10866_));
 sky130_fd_sc_hd__inv_16 _16320_ (.A(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_897 ();
 sky130_fd_sc_hd__mux2i_1 _16323_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10869_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10870_));
 sky130_fd_sc_hd__nand2_1 _16325_ (.A(net3948),
    .B(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__o21a_4 _16326_ (.A1(net3948),
    .A2(_10869_),
    .B1(_10871_),
    .X(_10872_));
 sky130_fd_sc_hd__clkinv_16 _16327_ (.A(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_895 ();
 sky130_fd_sc_hd__mux2i_1 _16330_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10875_));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10876_));
 sky130_fd_sc_hd__nand2_1 _16332_ (.A(net3948),
    .B(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__o21a_4 _16333_ (.A1(net3948),
    .A2(_10875_),
    .B1(_10877_),
    .X(_10878_));
 sky130_fd_sc_hd__clkinv_16 _16334_ (.A(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_893 ();
 sky130_fd_sc_hd__mux2i_1 _16337_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10881_));
 sky130_fd_sc_hd__mux2_4 _16338_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10882_));
 sky130_fd_sc_hd__nand2_1 _16339_ (.A(net3948),
    .B(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__o21a_4 _16340_ (.A1(net3948),
    .A2(_10881_),
    .B1(_10883_),
    .X(_10884_));
 sky130_fd_sc_hd__inv_8 _16341_ (.A(_10884_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[3] ));
 sky130_fd_sc_hd__mux2i_1 _16342_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10885_));
 sky130_fd_sc_hd__mux2_8 _16343_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10886_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(net3948),
    .B(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__o21a_4 _16345_ (.A1(net3948),
    .A2(_10885_),
    .B1(_10887_),
    .X(_10888_));
 sky130_fd_sc_hd__inv_4 _16346_ (.A(_10888_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[2] ));
 sky130_fd_sc_hd__mux2i_1 _16347_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10889_));
 sky130_fd_sc_hd__mux2_8 _16348_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10890_));
 sky130_fd_sc_hd__nand2_1 _16349_ (.A(net3948),
    .B(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__o21ai_4 _16350_ (.A1(net3948),
    .A2(_10889_),
    .B1(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_892 ();
 sky130_fd_sc_hd__mux2i_1 _16352_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10893_));
 sky130_fd_sc_hd__mux2_4 _16353_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10894_));
 sky130_fd_sc_hd__nand2_1 _16354_ (.A(net3948),
    .B(_10894_),
    .Y(_10895_));
 sky130_fd_sc_hd__o21a_4 _16355_ (.A1(net3948),
    .A2(_10893_),
    .B1(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_891 ();
 sky130_fd_sc_hd__clkinv_8 _16357_ (.A(_10896_),
    .Y(_10898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_890 ();
 sky130_fd_sc_hd__mux2_1 _16359_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_889 ();
 sky130_fd_sc_hd__mux2i_1 _16361_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10900_));
 sky130_fd_sc_hd__inv_1 _16362_ (.A(_10900_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ));
 sky130_fd_sc_hd__mux2i_1 _16363_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10901_));
 sky130_fd_sc_hd__inv_1 _16364_ (.A(_10901_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_888 ();
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ));
 sky130_fd_sc_hd__mux2_4 _16367_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ));
 sky130_fd_sc_hd__mux2i_1 _16369_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10903_));
 sky130_fd_sc_hd__inv_1 _16370_ (.A(_10903_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ));
 sky130_fd_sc_hd__mux2i_1 _16371_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10904_));
 sky130_fd_sc_hd__inv_1 _16372_ (.A(_10904_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ));
 sky130_fd_sc_hd__mux2_1 _16373_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ));
 sky130_fd_sc_hd__mux2i_1 _16374_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10905_));
 sky130_fd_sc_hd__inv_1 _16375_ (.A(_10905_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ));
 sky130_fd_sc_hd__mux2i_1 _16376_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10906_));
 sky130_fd_sc_hd__inv_1 _16377_ (.A(_10906_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ));
 sky130_fd_sc_hd__mux2i_1 _16378_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10907_));
 sky130_fd_sc_hd__inv_1 _16379_ (.A(_10907_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ));
 sky130_fd_sc_hd__mux2_1 _16380_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ));
 sky130_fd_sc_hd__mux2_1 _16381_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ));
 sky130_fd_sc_hd__mux2_1 _16382_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ));
 sky130_fd_sc_hd__o31ai_1 _16384_ (.A1(net60),
    .A2(core_busy_q),
    .A3(_10821_),
    .B1(fetch_enable_q),
    .Y(net150));
 sky130_fd_sc_hd__nand2b_1 _16385_ (.A_N(net149),
    .B(net150),
    .Y(_00008_));
 sky130_fd_sc_hd__clkinvlp_4 _16386_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_10908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_885 ();
 sky130_fd_sc_hd__nand2_4 _16390_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(net128),
    .Y(_10912_));
 sky130_fd_sc_hd__nor4_2 _16391_ (.A(_10908_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .D(_10912_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ));
 sky130_fd_sc_hd__inv_2 _16392_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10913_));
 sky130_fd_sc_hd__nor2_4 _16393_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .B(_10912_),
    .Y(_10914_));
 sky130_fd_sc_hd__and3_1 _16394_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .X(_10915_));
 sky130_fd_sc_hd__a31oi_1 _16395_ (.A1(_10913_),
    .A2(net104),
    .A3(net103),
    .B1(_10915_),
    .Y(_10916_));
 sky130_fd_sc_hd__mux2i_1 _16396_ (.A0(net94),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10917_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(_10916_),
    .B(_10917_),
    .Y(_10918_));
 sky130_fd_sc_hd__nand2_2 _16398_ (.A(net3948),
    .B(_10918_),
    .Y(_10919_));
 sky130_fd_sc_hd__nor2_1 _16399_ (.A(_10908_),
    .B(_10919_),
    .Y(_10920_));
 sky130_fd_sc_hd__a21oi_1 _16400_ (.A1(_10914_),
    .A2(_10919_),
    .B1(_10920_),
    .Y(_10921_));
 sky130_fd_sc_hd__nor3_1 _16401_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(_10914_),
    .C(_10919_),
    .Y(_10922_));
 sky130_fd_sc_hd__a211oi_4 _16402_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(net3785),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Y(_10923_));
 sky130_fd_sc_hd__nand2_8 _16403_ (.A(net3756),
    .B(_10923_),
    .Y(_10924_));
 sky130_fd_sc_hd__o21ai_0 _16404_ (.A1(\id_stage_i.id_fsm_q ),
    .A2(_10779_),
    .B1(_10924_),
    .Y(_10925_));
 sky130_fd_sc_hd__a21boi_0 _16405_ (.A1(\id_stage_i.id_fsm_q ),
    .A2(_10654_),
    .B1_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_10926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_884 ();
 sky130_fd_sc_hd__xor2_1 _16407_ (.A(_10393_),
    .B(net3587),
    .X(_10928_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_883 ();
 sky130_fd_sc_hd__o21a_4 _16409_ (.A1(net3939),
    .A2(_08093_),
    .B1(_08065_),
    .X(_10930_));
 sky130_fd_sc_hd__o221ai_4 _16410_ (.A1(_08063_),
    .A2(net394),
    .B1(_10930_),
    .B2(net3942),
    .C1(_08070_),
    .Y(_10931_));
 sky130_fd_sc_hd__and2_4 _16411_ (.A(_08087_),
    .B(_08092_),
    .X(_10932_));
 sky130_fd_sc_hd__nand2_1 _16412_ (.A(_08010_),
    .B(_08058_),
    .Y(_10933_));
 sky130_fd_sc_hd__nand2_1 _16413_ (.A(_08093_),
    .B(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__nor3_1 _16414_ (.A(_08019_),
    .B(_08014_),
    .C(_08093_),
    .Y(_10935_));
 sky130_fd_sc_hd__a21oi_2 _16415_ (.A1(net3940),
    .A2(_10934_),
    .B1(_10935_),
    .Y(_10936_));
 sky130_fd_sc_hd__and3_4 _16416_ (.A(_10932_),
    .B(net3725),
    .C(_10936_),
    .X(_10937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_882 ();
 sky130_fd_sc_hd__nand2_2 _16418_ (.A(_10931_),
    .B(_10937_),
    .Y(_10939_));
 sky130_fd_sc_hd__clkinv_2 _16419_ (.A(_10931_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(net384),
    .B(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__and2_4 _16421_ (.A(_10932_),
    .B(_10936_),
    .X(_10942_));
 sky130_fd_sc_hd__o221a_1 _16422_ (.A1(net383),
    .A2(_10939_),
    .B1(_10941_),
    .B2(_10942_),
    .C1(_08088_),
    .X(_10943_));
 sky130_fd_sc_hd__o21ai_2 _16423_ (.A1(_08051_),
    .A2(_10943_),
    .B1(_10932_),
    .Y(_10944_));
 sky130_fd_sc_hd__or2_4 _16424_ (.A(net384),
    .B(_10931_),
    .X(_10945_));
 sky130_fd_sc_hd__nand2_2 _16425_ (.A(net384),
    .B(_10931_),
    .Y(_10946_));
 sky130_fd_sc_hd__nand2_4 _16426_ (.A(_08088_),
    .B(_08032_),
    .Y(_10947_));
 sky130_fd_sc_hd__a21oi_4 _16427_ (.A1(_10945_),
    .A2(_10946_),
    .B1(_10947_),
    .Y(_10948_));
 sky130_fd_sc_hd__mux2_1 _16428_ (.A0(_10944_),
    .A1(_10948_),
    .S(net3470),
    .X(_10949_));
 sky130_fd_sc_hd__o221ai_1 _16429_ (.A1(_08093_),
    .A2(_10936_),
    .B1(_10947_),
    .B2(net3725),
    .C1(_10932_),
    .Y(_10950_));
 sky130_fd_sc_hd__a32oi_1 _16430_ (.A1(_08088_),
    .A2(_08032_),
    .A3(_10937_),
    .B1(_10950_),
    .B2(net383),
    .Y(_10951_));
 sky130_fd_sc_hd__nor2_2 _16431_ (.A(_10940_),
    .B(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__mux2i_1 _16432_ (.A0(_10944_),
    .A1(_10948_),
    .S(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__nand3b_1 _16433_ (.A_N(net3587),
    .B(_10953_),
    .C(_10393_),
    .Y(_10954_));
 sky130_fd_sc_hd__xnor2_1 _16434_ (.A(_10952_),
    .B(_10948_),
    .Y(_10955_));
 sky130_fd_sc_hd__nand3b_1 _16435_ (.A_N(_10393_),
    .B(net3587),
    .C(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__o211ai_1 _16436_ (.A1(_10928_),
    .A2(_10949_),
    .B1(_10954_),
    .C1(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__nor3_1 _16437_ (.A(net3725),
    .B(_10941_),
    .C(_10947_),
    .Y(_10958_));
 sky130_fd_sc_hd__nor3_1 _16438_ (.A(_10944_),
    .B(_10948_),
    .C(_10958_),
    .Y(_10959_));
 sky130_fd_sc_hd__mux2i_1 _16439_ (.A0(_10958_),
    .A1(_10959_),
    .S(_10736_),
    .Y(_10960_));
 sky130_fd_sc_hd__a2111oi_2 _16440_ (.A1(net3462),
    .A2(net3461),
    .B1(_07874_),
    .C1(_07884_),
    .D1(_10780_),
    .Y(\id_stage_i.branch_set_d ));
 sky130_fd_sc_hd__a221o_4 _16441_ (.A1(_10542_),
    .A2(_10925_),
    .B1(_10926_),
    .B2(_10657_),
    .C1(\id_stage_i.branch_set_d ),
    .X(_10961_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_881 ();
 sky130_fd_sc_hd__nand3b_1 _16443_ (.A_N(net3933),
    .B(net3775),
    .C(net3781),
    .Y(_10963_));
 sky130_fd_sc_hd__and3_4 _16444_ (.A(net3940),
    .B(net3750),
    .C(_10963_),
    .X(_10964_));
 sky130_fd_sc_hd__nand2_8 _16445_ (.A(net3943),
    .B(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__nor3_1 _16446_ (.A(net3895),
    .B(net3858),
    .C(_10512_),
    .Y(_10966_));
 sky130_fd_sc_hd__nor3_1 _16447_ (.A(net3851),
    .B(_10508_),
    .C(_10965_),
    .Y(_10967_));
 sky130_fd_sc_hd__a21oi_1 _16448_ (.A1(_10965_),
    .A2(_10966_),
    .B1(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__nand3_1 _16449_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(net3839),
    .C(_10502_),
    .Y(_10969_));
 sky130_fd_sc_hd__or3_4 _16450_ (.A(_10546_),
    .B(_10968_),
    .C(_10969_),
    .X(_10970_));
 sky130_fd_sc_hd__nand2b_1 _16451_ (.A_N(_10504_),
    .B(_10516_),
    .Y(_10971_));
 sky130_fd_sc_hd__and3_4 _16452_ (.A(_10655_),
    .B(_10970_),
    .C(_10971_),
    .X(_10972_));
 sky130_fd_sc_hd__nand2b_1 _16453_ (.A_N(_10649_),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__a21oi_1 _16454_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(\cs_registers_i.dcsr_q[2] ),
    .B1(net60),
    .Y(_10974_));
 sky130_fd_sc_hd__nor2_2 _16455_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__a211oi_1 _16456_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_10973_),
    .B1(_10975_),
    .C1(_10823_),
    .Y(_10976_));
 sky130_fd_sc_hd__clkinv_1 _16457_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_10977_));
 sky130_fd_sc_hd__nand2_4 _16458_ (.A(_10977_),
    .B(_10498_),
    .Y(_10978_));
 sky130_fd_sc_hd__o311ai_2 _16459_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_10538_),
    .A3(_10976_),
    .B1(_10978_),
    .C1(_10500_),
    .Y(_10979_));
 sky130_fd_sc_hd__a2111oi_2 _16460_ (.A1(_10913_),
    .A2(_10921_),
    .B1(_10922_),
    .C1(_10961_),
    .D1(_10979_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux2_1 _16461_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_10738_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .S(_10738_),
    .X(_00011_));
 sky130_fd_sc_hd__and3_4 _16463_ (.A(net3612),
    .B(net3673),
    .C(_10690_),
    .X(_10980_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_880 ();
 sky130_fd_sc_hd__nand2_1 _16465_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_10980_),
    .Y(_10982_));
 sky130_fd_sc_hd__o21ai_0 _16466_ (.A1(_08169_),
    .A2(_10683_),
    .B1(_10982_),
    .Y(_00012_));
 sky130_fd_sc_hd__nand2_1 _16467_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_10679_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand2_8 _16468_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(_10683_),
    .Y(_10984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_879 ();
 sky130_fd_sc_hd__nand2_1 _16470_ (.A(_10983_),
    .B(_10984_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(_10980_),
    .Y(_10986_));
 sky130_fd_sc_hd__o21ai_0 _16472_ (.A1(_10686_),
    .A2(_10683_),
    .B1(_10986_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_2 _16473_ (.A(net3614),
    .B(_10571_),
    .Y(_10987_));
 sky130_fd_sc_hd__nor4_4 _16474_ (.A(_10546_),
    .B(_10627_),
    .C(_10636_),
    .D(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_878 ();
 sky130_fd_sc_hd__nand2_2 _16476_ (.A(net3551),
    .B(net3501),
    .Y(_10990_));
 sky130_fd_sc_hd__nand3_4 _16477_ (.A(net3940),
    .B(net3750),
    .C(_10963_),
    .Y(_10991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_877 ();
 sky130_fd_sc_hd__nand2_8 _16479_ (.A(_10557_),
    .B(_10596_),
    .Y(_10993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_875 ();
 sky130_fd_sc_hd__nor2_4 _16482_ (.A(_10549_),
    .B(_10600_),
    .Y(_10996_));
 sky130_fd_sc_hd__nand4_1 _16483_ (.A(net3618),
    .B(net3616),
    .C(net3614),
    .D(_10557_),
    .Y(_10997_));
 sky130_fd_sc_hd__nand2b_4 _16484_ (.A_N(_10997_),
    .B(net353),
    .Y(_10998_));
 sky130_fd_sc_hd__nor2b_4 _16485_ (.A(_10998_),
    .B_N(net3625),
    .Y(_10999_));
 sky130_fd_sc_hd__nor2_4 _16486_ (.A(_10570_),
    .B(_10597_),
    .Y(_11000_));
 sky130_fd_sc_hd__nor3_4 _16487_ (.A(net3625),
    .B(_10997_),
    .C(_10577_),
    .Y(_11001_));
 sky130_fd_sc_hd__and2_4 _16488_ (.A(_10572_),
    .B(_11001_),
    .X(_11002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_874 ();
 sky130_fd_sc_hd__and2_4 _16490_ (.A(_11001_),
    .B(_10580_),
    .X(_11004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_873 ();
 sky130_fd_sc_hd__a222oi_1 _16492_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11002_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .C2(_11004_),
    .Y(_11006_));
 sky130_fd_sc_hd__a22oi_2 _16493_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(_11002_),
    .B1(_11004_),
    .B2(\cs_registers_i.mhpmcounter[1888] ),
    .Y(_11007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_872 ();
 sky130_fd_sc_hd__nand2_8 _16495_ (.A(net3621),
    .B(_10616_),
    .Y(_11009_));
 sky130_fd_sc_hd__o22ai_4 _16496_ (.A1(_10996_),
    .A2(_11006_),
    .B1(_11007_),
    .B2(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_871 ();
 sky130_fd_sc_hd__nor3_4 _16498_ (.A(net3619),
    .B(net3595),
    .C(_10566_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand2_1 _16499_ (.A(_10592_),
    .B(_11012_),
    .Y(_11013_));
 sky130_fd_sc_hd__nand2_2 _16500_ (.A(_10557_),
    .B(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__and3_4 _16501_ (.A(net3586),
    .B(_11014_),
    .C(_10999_),
    .X(_11015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_870 ();
 sky130_fd_sc_hd__nand3_2 _16503_ (.A(net3618),
    .B(net3616),
    .C(_10557_),
    .Y(_11017_));
 sky130_fd_sc_hd__or3_4 _16504_ (.A(net3586),
    .B(net3614),
    .C(_11017_),
    .X(_11018_));
 sky130_fd_sc_hd__or4_4 _16505_ (.A(_10552_),
    .B(_10556_),
    .C(_10560_),
    .D(_11018_),
    .X(_11019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_868 ();
 sky130_fd_sc_hd__nand2_4 _16508_ (.A(net3619),
    .B(_10616_),
    .Y(_11022_));
 sky130_fd_sc_hd__nor2_4 _16509_ (.A(_11019_),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__nor2_4 _16510_ (.A(_11019_),
    .B(_11009_),
    .Y(_11024_));
 sky130_fd_sc_hd__a222oi_1 _16511_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11015_),
    .B1(_11023_),
    .B2(\cs_registers_i.dscratch1_q[0] ),
    .C1(_11024_),
    .C2(\cs_registers_i.dscratch0_q[0] ),
    .Y(_11025_));
 sky130_fd_sc_hd__or3_4 _16512_ (.A(_08779_),
    .B(_10998_),
    .C(_10587_),
    .X(_11026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_867 ();
 sky130_fd_sc_hd__nor2_4 _16514_ (.A(_10585_),
    .B(_11026_),
    .Y(_11028_));
 sky130_fd_sc_hd__nor2_4 _16515_ (.A(_11026_),
    .B(_10618_),
    .Y(_11029_));
 sky130_fd_sc_hd__nor4_4 _16516_ (.A(_10556_),
    .B(_10560_),
    .C(_11018_),
    .D(_10585_),
    .Y(_11030_));
 sky130_fd_sc_hd__a222oi_1 _16517_ (.A1(\cs_registers_i.mscratch_q[0] ),
    .A2(_11028_),
    .B1(_11029_),
    .B2(\cs_registers_i.mtval_q[0] ),
    .C1(\cs_registers_i.dcsr_q[0] ),
    .C2(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__nor3_4 _16518_ (.A(net3625),
    .B(_11018_),
    .C(_10603_),
    .Y(_11032_));
 sky130_fd_sc_hd__nor2_2 _16519_ (.A(_11026_),
    .B(_10612_),
    .Y(_11033_));
 sky130_fd_sc_hd__a22oi_1 _16520_ (.A1(net62),
    .A2(_11032_),
    .B1(_11033_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .Y(_11034_));
 sky130_fd_sc_hd__nor2_4 _16521_ (.A(_10576_),
    .B(_11026_),
    .Y(_11035_));
 sky130_fd_sc_hd__or2_4 _16522_ (.A(_10998_),
    .B(_10593_),
    .X(_11036_));
 sky130_fd_sc_hd__nor2_4 _16523_ (.A(_11036_),
    .B(_10614_),
    .Y(_11037_));
 sky130_fd_sc_hd__a21oi_1 _16524_ (.A1(\cs_registers_i.csr_mepc_o[0] ),
    .A2(_11035_),
    .B1(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand4_1 _16525_ (.A(_11025_),
    .B(_11031_),
    .C(_11034_),
    .D(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__a21oi_4 _16526_ (.A1(_10993_),
    .A2(_11010_),
    .B1(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__o21ai_1 _16527_ (.A1(_10991_),
    .A2(_11040_),
    .B1(net3620),
    .Y(_11041_));
 sky130_fd_sc_hd__o21ai_4 _16528_ (.A1(net3620),
    .A2(_10965_),
    .B1(_11041_),
    .Y(_11042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_865 ();
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_10990_),
    .Y(_11045_));
 sky130_fd_sc_hd__o21ai_0 _16532_ (.A1(_10990_),
    .A2(_11042_),
    .B1(_11045_),
    .Y(_00015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_863 ();
 sky130_fd_sc_hd__a22oi_2 _16535_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A2(_10579_),
    .B1(_10581_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .Y(_11048_));
 sky130_fd_sc_hd__and2_4 _16536_ (.A(net3625),
    .B(_10589_),
    .X(_11049_));
 sky130_fd_sc_hd__a222oi_1 _16537_ (.A1(\cs_registers_i.mhpmcounter[1858] ),
    .A2(_10579_),
    .B1(_10581_),
    .B2(\cs_registers_i.mhpmcounter[1890] ),
    .C1(_11049_),
    .C2(_11000_),
    .Y(_11050_));
 sky130_fd_sc_hd__o22ai_4 _16538_ (.A1(_10996_),
    .A2(_11048_),
    .B1(_11050_),
    .B2(_11009_),
    .Y(_11051_));
 sky130_fd_sc_hd__and3_4 _16539_ (.A(net3586),
    .B(_11014_),
    .C(_11049_),
    .X(_11052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_861 ();
 sky130_fd_sc_hd__or4_4 _16542_ (.A(net3586),
    .B(_10556_),
    .C(_10560_),
    .D(_10564_),
    .X(_11055_));
 sky130_fd_sc_hd__nand2b_4 _16543_ (.A_N(_11055_),
    .B(_10567_),
    .Y(_11056_));
 sky130_fd_sc_hd__nor2_4 _16544_ (.A(_11009_),
    .B(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_860 ();
 sky130_fd_sc_hd__nor2_4 _16546_ (.A(_11022_),
    .B(_11056_),
    .Y(_11059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_859 ();
 sky130_fd_sc_hd__a222oi_1 _16548_ (.A1(\cs_registers_i.mcountinhibit_q[2] ),
    .A2(_11052_),
    .B1(_11057_),
    .B2(\cs_registers_i.dscratch0_q[2] ),
    .C1(_11059_),
    .C2(\cs_registers_i.dscratch1_q[2] ),
    .Y(_11061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_858 ();
 sky130_fd_sc_hd__nor2_4 _16550_ (.A(_10585_),
    .B(_11055_),
    .Y(_11063_));
 sky130_fd_sc_hd__a22oi_2 _16551_ (.A1(\cs_registers_i.mscratch_q[2] ),
    .A2(net3540),
    .B1(_11063_),
    .B2(\cs_registers_i.dcsr_q[2] ),
    .Y(_11064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_857 ();
 sky130_fd_sc_hd__a22oi_2 _16553_ (.A1(\cs_registers_i.mcause_q[2] ),
    .A2(_10613_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[2] ),
    .Y(_11066_));
 sky130_fd_sc_hd__nand3_4 _16554_ (.A(_10557_),
    .B(_10600_),
    .C(_10601_),
    .Y(_11067_));
 sky130_fd_sc_hd__nor3_1 _16555_ (.A(net3625),
    .B(net3586),
    .C(_10564_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand2_2 _16556_ (.A(_10572_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__nor2_4 _16557_ (.A(_11067_),
    .B(_11069_),
    .Y(_11070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_855 ();
 sky130_fd_sc_hd__inv_6 _16560_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .Y(_11073_));
 sky130_fd_sc_hd__o21ai_2 _16561_ (.A1(_11073_),
    .A2(_10590_),
    .B1(_10594_),
    .Y(_11074_));
 sky130_fd_sc_hd__inv_1 _16562_ (.A(_10576_),
    .Y(_11075_));
 sky130_fd_sc_hd__nor2_4 _16563_ (.A(_10576_),
    .B(_11055_),
    .Y(_11076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_854 ();
 sky130_fd_sc_hd__a222oi_1 _16565_ (.A1(net84),
    .A2(_11070_),
    .B1(_11074_),
    .B2(_11075_),
    .C1(_11076_),
    .C2(\cs_registers_i.csr_depc_o[2] ),
    .Y(_11078_));
 sky130_fd_sc_hd__nand4_1 _16566_ (.A(_11061_),
    .B(_11064_),
    .C(_11066_),
    .D(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__a21oi_4 _16567_ (.A1(_10993_),
    .A2(_11051_),
    .B1(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__o21ai_1 _16568_ (.A1(_10991_),
    .A2(_11080_),
    .B1(net3598),
    .Y(_11081_));
 sky130_fd_sc_hd__o21ai_4 _16569_ (.A1(net3598),
    .A2(_10965_),
    .B1(_11081_),
    .Y(_11082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_853 ();
 sky130_fd_sc_hd__nand2_1 _16571_ (.A(\cs_registers_i.mcountinhibit_q[2] ),
    .B(_10990_),
    .Y(_11084_));
 sky130_fd_sc_hd__o21ai_0 _16572_ (.A1(_10990_),
    .A2(_11082_),
    .B1(_11084_),
    .Y(_00016_));
 sky130_fd_sc_hd__o21ai_4 _16573_ (.A1(_08737_),
    .A2(_10566_),
    .B1(_10557_),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_4 _16574_ (.A(_11085_),
    .B(_10988_),
    .Y(_11086_));
 sky130_fd_sc_hd__or3_4 _16575_ (.A(_10996_),
    .B(_10583_),
    .C(_11086_),
    .X(_11087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_852 ();
 sky130_fd_sc_hd__nand2_8 _16577_ (.A(_10580_),
    .B(_10578_),
    .Y(_11089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_851 ();
 sky130_fd_sc_hd__nor2_4 _16579_ (.A(_11089_),
    .B(_11087_),
    .Y(_11091_));
 sky130_fd_sc_hd__a21oi_1 _16580_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11087_),
    .B1(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__a21oi_4 _16581_ (.A1(net3586),
    .A2(_10551_),
    .B1(_10549_),
    .Y(_11093_));
 sky130_fd_sc_hd__nand2_2 _16582_ (.A(_08779_),
    .B(_10563_),
    .Y(_11094_));
 sky130_fd_sc_hd__nand3_1 _16583_ (.A(net3618),
    .B(net3616),
    .C(_10557_),
    .Y(_11095_));
 sky130_fd_sc_hd__nor4_1 _16584_ (.A(_10587_),
    .B(_10616_),
    .C(_11094_),
    .D(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_850 ();
 sky130_fd_sc_hd__nor2_4 _16586_ (.A(_10594_),
    .B(_11067_),
    .Y(_11098_));
 sky130_fd_sc_hd__a2111oi_0 _16587_ (.A1(_10622_),
    .A2(_11096_),
    .B1(net3550),
    .C1(_11098_),
    .D1(_10613_),
    .Y(_11099_));
 sky130_fd_sc_hd__nand2_1 _16588_ (.A(net3625),
    .B(_10589_),
    .Y(_11100_));
 sky130_fd_sc_hd__o21ai_0 _16589_ (.A1(_10554_),
    .A2(_11100_),
    .B1(_11056_),
    .Y(_11101_));
 sky130_fd_sc_hd__or2_4 _16590_ (.A(_10606_),
    .B(_11052_),
    .X(_11102_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(_11000_),
    .B(_11049_),
    .Y(_11103_));
 sky130_fd_sc_hd__nor2_4 _16592_ (.A(_10590_),
    .B(_11067_),
    .Y(_11104_));
 sky130_fd_sc_hd__nor2_1 _16593_ (.A(_11070_),
    .B(_11104_),
    .Y(_11105_));
 sky130_fd_sc_hd__nor4_1 _16594_ (.A(net3540),
    .B(_10625_),
    .C(_10595_),
    .D(net3539),
    .Y(_11106_));
 sky130_fd_sc_hd__nand3_1 _16595_ (.A(_11103_),
    .B(_11105_),
    .C(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__a211oi_1 _16596_ (.A1(_10553_),
    .A2(_11101_),
    .B1(_11102_),
    .C1(_11107_),
    .Y(_11108_));
 sky130_fd_sc_hd__nand3_1 _16597_ (.A(_10583_),
    .B(_11099_),
    .C(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__nor2_2 _16598_ (.A(_10546_),
    .B(_10987_),
    .Y(_11110_));
 sky130_fd_sc_hd__o2111ai_2 _16599_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_11056_),
    .B1(_11109_),
    .C1(_11110_),
    .D1(_10635_),
    .Y(_11111_));
 sky130_fd_sc_hd__nor4_4 _16600_ (.A(_10996_),
    .B(_11093_),
    .C(_10583_),
    .D(_11111_),
    .Y(_11112_));
 sky130_fd_sc_hd__nor2_4 _16601_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_849 ();
 sky130_fd_sc_hd__nor2_4 _16603_ (.A(_10581_),
    .B(_11087_),
    .Y(_11115_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_848 ();
 sky130_fd_sc_hd__a22oi_1 _16605_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_11113_),
    .B1(_11115_),
    .B2(_11042_),
    .Y(_11117_));
 sky130_fd_sc_hd__o21a_1 _16606_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_11092_),
    .B1(_11117_),
    .X(_00017_));
 sky130_fd_sc_hd__or4_4 _16607_ (.A(_10996_),
    .B(_11093_),
    .C(_10583_),
    .D(_11111_),
    .X(_11118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_847 ();
 sky130_fd_sc_hd__nor2_4 _16609_ (.A(_10581_),
    .B(_11118_),
    .Y(_11120_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_843 ();
 sky130_fd_sc_hd__a21oi_1 _16614_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(net3539),
    .B1(_11052_),
    .Y(_11125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_842 ();
 sky130_fd_sc_hd__a22oi_2 _16616_ (.A1(net63),
    .A2(net3546),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[10] ),
    .Y(_11127_));
 sky130_fd_sc_hd__nand2_4 _16617_ (.A(_11125_),
    .B(_11127_),
    .Y(_11128_));
 sky130_fd_sc_hd__a221oi_1 _16618_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[10] ),
    .C1(_11128_),
    .Y(_11129_));
 sky130_fd_sc_hd__nand2_8 _16619_ (.A(_10572_),
    .B(_10578_),
    .Y(_11130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_836 ();
 sky130_fd_sc_hd__a22oi_2 _16626_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1866] ),
    .Y(_11137_));
 sky130_fd_sc_hd__a22oi_2 _16627_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1898] ),
    .Y(_11138_));
 sky130_fd_sc_hd__o22ai_4 _16628_ (.A1(_11130_),
    .A2(_11137_),
    .B1(_11138_),
    .B2(_11089_),
    .Y(_11139_));
 sky130_fd_sc_hd__nand2_2 _16629_ (.A(_10993_),
    .B(_11139_),
    .Y(_11140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_835 ();
 sky130_fd_sc_hd__a222oi_1 _16631_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[10] ),
    .C1(net3566),
    .C2(\cs_registers_i.csr_depc_o[10] ),
    .Y(_11142_));
 sky130_fd_sc_hd__and3_4 _16632_ (.A(_11129_),
    .B(_11140_),
    .C(net3528),
    .X(_11143_));
 sky130_fd_sc_hd__nor3_1 _16633_ (.A(net3592),
    .B(_10991_),
    .C(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__a21oi_4 _16634_ (.A1(net3592),
    .A2(_10965_),
    .B1(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_834 ();
 sky130_fd_sc_hd__nor3_4 _16636_ (.A(_10996_),
    .B(_10583_),
    .C(_11086_),
    .Y(_11147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_833 ();
 sky130_fd_sc_hd__nand2_4 _16638_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .Y(_11149_));
 sky130_fd_sc_hd__and3_4 _16639_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .X(_11150_));
 sky130_fd_sc_hd__nand3_4 _16640_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .C(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__nor3_4 _16641_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11149_),
    .C(_11151_),
    .Y(_11152_));
 sky130_fd_sc_hd__nand3_1 _16642_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .C(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(net3484),
    .B(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__a211oi_1 _16644_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(_11154_),
    .B1(_11115_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .Y(_11155_));
 sky130_fd_sc_hd__nand4_1 _16645_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .D(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .Y(_11156_));
 sky130_fd_sc_hd__nor2_4 _16646_ (.A(_11149_),
    .B(_11151_),
    .Y(_11157_));
 sky130_fd_sc_hd__nor4b_2 _16647_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11156_),
    .C(net3484),
    .D_N(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__a211oi_1 _16648_ (.A1(_11120_),
    .A2(_11145_),
    .B1(_11155_),
    .C1(_11158_),
    .Y(_00018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_832 ();
 sky130_fd_sc_hd__a22oi_2 _16650_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1867] ),
    .Y(_11160_));
 sky130_fd_sc_hd__a22oi_2 _16651_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1899] ),
    .Y(_11161_));
 sky130_fd_sc_hd__o22ai_4 _16652_ (.A1(_11130_),
    .A2(_11160_),
    .B1(_11161_),
    .B2(_11089_),
    .Y(_11162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_830 ();
 sky130_fd_sc_hd__a222oi_1 _16655_ (.A1(net129),
    .A2(_11104_),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[11] ),
    .C1(_11063_),
    .C2(\cs_registers_i.dcsr_q[11] ),
    .Y(_11165_));
 sky130_fd_sc_hd__a22oi_2 _16656_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(net3550),
    .B1(net3546),
    .B2(net64),
    .Y(_11166_));
 sky130_fd_sc_hd__a21oi_2 _16657_ (.A1(\cs_registers_i.mstatus_q[2] ),
    .A2(_10595_),
    .B1(_11052_),
    .Y(_11167_));
 sky130_fd_sc_hd__nand3_4 _16658_ (.A(_11165_),
    .B(_11166_),
    .C(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__a22oi_2 _16659_ (.A1(\cs_registers_i.mtval_q[11] ),
    .A2(net3539),
    .B1(_11076_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .Y(_11169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_828 ();
 sky130_fd_sc_hd__a22oi_2 _16662_ (.A1(\cs_registers_i.mie_q[15] ),
    .A2(_11098_),
    .B1(_10625_),
    .B2(\cs_registers_i.csr_mepc_o[11] ),
    .Y(_11172_));
 sky130_fd_sc_hd__a22oi_2 _16663_ (.A1(\cs_registers_i.dscratch0_q[11] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[11] ),
    .Y(_11173_));
 sky130_fd_sc_hd__nand3_4 _16664_ (.A(_11169_),
    .B(_11172_),
    .C(_11173_),
    .Y(_11174_));
 sky130_fd_sc_hd__a211oi_4 _16665_ (.A1(_10993_),
    .A2(_11162_),
    .B1(_11168_),
    .C1(_11174_),
    .Y(_11175_));
 sky130_fd_sc_hd__nor3_1 _16666_ (.A(_08988_),
    .B(_10991_),
    .C(_11175_),
    .Y(_11176_));
 sky130_fd_sc_hd__a21oi_4 _16667_ (.A1(_08988_),
    .A2(_10965_),
    .B1(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_827 ();
 sky130_fd_sc_hd__and2_0 _16669_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .B(_11158_),
    .X(_11179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_826 ();
 sky130_fd_sc_hd__nor3_1 _16671_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .B(_11120_),
    .C(_11158_),
    .Y(_11181_));
 sky130_fd_sc_hd__a211oi_1 _16672_ (.A1(_11115_),
    .A2(_11177_),
    .B1(_11179_),
    .C1(_11181_),
    .Y(_00019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_822 ();
 sky130_fd_sc_hd__a22oi_2 _16677_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1900] ),
    .Y(_11186_));
 sky130_fd_sc_hd__a22oi_1 _16678_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1868] ),
    .Y(_11187_));
 sky130_fd_sc_hd__o22ai_4 _16679_ (.A1(_11089_),
    .A2(_11186_),
    .B1(_11187_),
    .B2(_11130_),
    .Y(_11188_));
 sky130_fd_sc_hd__a22o_1 _16680_ (.A1(\cs_registers_i.csr_mtvec_o[12] ),
    .A2(net3550),
    .B1(_10595_),
    .B2(\cs_registers_i.mstatus_q[3] ),
    .X(_11189_));
 sky130_fd_sc_hd__a221oi_2 _16681_ (.A1(\cs_registers_i.mtval_q[12] ),
    .A2(net3539),
    .B1(_11063_),
    .B2(\cs_registers_i.dcsr_q[12] ),
    .C1(_11189_),
    .Y(_11190_));
 sky130_fd_sc_hd__a22oi_2 _16682_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(net3538),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .Y(_11191_));
 sky130_fd_sc_hd__a22oi_2 _16683_ (.A1(net65),
    .A2(net3546),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[12] ),
    .Y(_11192_));
 sky130_fd_sc_hd__nand3_4 _16684_ (.A(_11190_),
    .B(_11191_),
    .C(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__a221o_4 _16685_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[12] ),
    .C1(_11102_),
    .X(_11194_));
 sky130_fd_sc_hd__a211oi_4 _16686_ (.A1(_10993_),
    .A2(_11188_),
    .B1(_11193_),
    .C1(_11194_),
    .Y(_11195_));
 sky130_fd_sc_hd__nor3_1 _16687_ (.A(_09214_),
    .B(_10991_),
    .C(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__a21oi_4 _16688_ (.A1(_09214_),
    .A2(_10965_),
    .B1(_11196_),
    .Y(_11197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_821 ();
 sky130_fd_sc_hd__nor4bb_1 _16690_ (.A(_11112_),
    .B(_11156_),
    .C_N(_11152_),
    .D_N(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .Y(_11199_));
 sky130_fd_sc_hd__nand2_1 _16691_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .B(_11179_),
    .Y(_11200_));
 sky130_fd_sc_hd__o31ai_1 _16692_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_11120_),
    .A3(_11199_),
    .B1(_11200_),
    .Y(_11201_));
 sky130_fd_sc_hd__a21oi_1 _16693_ (.A1(_11115_),
    .A2(_11197_),
    .B1(_11201_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand2_4 _16694_ (.A(_11089_),
    .B(net3484),
    .Y(_11202_));
 sky130_fd_sc_hd__a22oi_2 _16695_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1901] ),
    .Y(_11203_));
 sky130_fd_sc_hd__a22oi_1 _16696_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1869] ),
    .Y(_11204_));
 sky130_fd_sc_hd__o22ai_4 _16697_ (.A1(_11089_),
    .A2(_11203_),
    .B1(_11204_),
    .B2(_11130_),
    .Y(_11205_));
 sky130_fd_sc_hd__a22o_1 _16698_ (.A1(net66),
    .A2(_11070_),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[13] ),
    .X(_11206_));
 sky130_fd_sc_hd__a221o_4 _16699_ (.A1(\cs_registers_i.mscratch_q[13] ),
    .A2(net3540),
    .B1(_11063_),
    .B2(\cs_registers_i.dcsr_q[13] ),
    .C1(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__a21oi_1 _16700_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(net3539),
    .B1(_11052_),
    .Y(_11208_));
 sky130_fd_sc_hd__a22oi_2 _16701_ (.A1(\cs_registers_i.csr_mtvec_o[13] ),
    .A2(net3550),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .Y(_11209_));
 sky130_fd_sc_hd__a22oi_1 _16702_ (.A1(\cs_registers_i.dscratch0_q[13] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[13] ),
    .Y(_11210_));
 sky130_fd_sc_hd__nand3_2 _16703_ (.A(_11208_),
    .B(_11209_),
    .C(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__a211oi_4 _16704_ (.A1(_10993_),
    .A2(_11205_),
    .B1(_11207_),
    .C1(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__nor3_1 _16705_ (.A(net3591),
    .B(_10991_),
    .C(_11212_),
    .Y(_11213_));
 sky130_fd_sc_hd__a21oi_4 _16706_ (.A1(net3591),
    .A2(_10965_),
    .B1(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_820 ();
 sky130_fd_sc_hd__nand2_2 _16708_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .Y(_11216_));
 sky130_fd_sc_hd__nor2_4 _16709_ (.A(_11156_),
    .B(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__a21oi_1 _16710_ (.A1(_11152_),
    .A2(_11217_),
    .B1(net3484),
    .Y(_11218_));
 sky130_fd_sc_hd__o21ai_0 _16711_ (.A1(_11091_),
    .A2(_11218_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .Y(_11219_));
 sky130_fd_sc_hd__nand4b_1 _16712_ (.A_N(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .B(_11087_),
    .C(_11152_),
    .D(_11217_),
    .Y(_11220_));
 sky130_fd_sc_hd__o211ai_1 _16713_ (.A1(_11202_),
    .A2(_11214_),
    .B1(_11219_),
    .C1(_11220_),
    .Y(_00021_));
 sky130_fd_sc_hd__nor2_4 _16714_ (.A(_10576_),
    .B(_10565_),
    .Y(_11221_));
 sky130_fd_sc_hd__a222oi_1 _16715_ (.A1(\cs_registers_i.csr_mtvec_o[14] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[14] ),
    .C1(_11221_),
    .C2(\cs_registers_i.csr_depc_o[14] ),
    .Y(_11222_));
 sky130_fd_sc_hd__a22oi_1 _16716_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1902] ),
    .Y(_11223_));
 sky130_fd_sc_hd__a22oi_1 _16717_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1870] ),
    .Y(_11224_));
 sky130_fd_sc_hd__o22ai_2 _16718_ (.A1(_11089_),
    .A2(_11223_),
    .B1(_11224_),
    .B2(_11130_),
    .Y(_11225_));
 sky130_fd_sc_hd__nand2_2 _16719_ (.A(_11085_),
    .B(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__nor2_4 _16720_ (.A(_11022_),
    .B(_10568_),
    .Y(_11227_));
 sky130_fd_sc_hd__nor2_4 _16721_ (.A(_11009_),
    .B(_10568_),
    .Y(_11228_));
 sky130_fd_sc_hd__a21oi_1 _16722_ (.A1(\cs_registers_i.csr_mepc_o[14] ),
    .A2(net3538),
    .B1(net3551),
    .Y(_11229_));
 sky130_fd_sc_hd__a22oi_1 _16723_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(net3539),
    .B1(net3552),
    .B2(net67),
    .Y(_11230_));
 sky130_fd_sc_hd__nand2_2 _16724_ (.A(_11229_),
    .B(_11230_),
    .Y(_11231_));
 sky130_fd_sc_hd__a221oi_1 _16725_ (.A1(\cs_registers_i.dscratch1_q[14] ),
    .A2(_11227_),
    .B1(_11228_),
    .B2(\cs_registers_i.dscratch0_q[14] ),
    .C1(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__and3_4 _16726_ (.A(net3527),
    .B(_11226_),
    .C(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__nor3_1 _16727_ (.A(net3589),
    .B(_10991_),
    .C(_11233_),
    .Y(_11234_));
 sky130_fd_sc_hd__a21oi_4 _16728_ (.A1(net3589),
    .A2(_10965_),
    .B1(_11234_),
    .Y(_11235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_819 ();
 sky130_fd_sc_hd__and4b_1 _16730_ (.A_N(\cs_registers_i.mcountinhibit_q[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .C(_11157_),
    .D(_11217_),
    .X(_11237_));
 sky130_fd_sc_hd__nand2_1 _16731_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .B(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_11112_),
    .B(_11238_),
    .Y(_11239_));
 sky130_fd_sc_hd__nand2_8 _16733_ (.A(_10581_),
    .B(net3484),
    .Y(_11240_));
 sky130_fd_sc_hd__nand3_1 _16734_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .B(_11157_),
    .C(_11217_),
    .Y(_11241_));
 sky130_fd_sc_hd__o21ai_0 _16735_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11241_),
    .B1(_11087_),
    .Y(_11242_));
 sky130_fd_sc_hd__a21oi_1 _16736_ (.A1(_11240_),
    .A2(_11242_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .Y(_11243_));
 sky130_fd_sc_hd__a211oi_1 _16737_ (.A1(_11120_),
    .A2(_11235_),
    .B1(_11239_),
    .C1(_11243_),
    .Y(_00022_));
 sky130_fd_sc_hd__a22oi_2 _16738_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1903] ),
    .Y(_11244_));
 sky130_fd_sc_hd__a22oi_1 _16739_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1871] ),
    .Y(_11245_));
 sky130_fd_sc_hd__o22ai_4 _16740_ (.A1(_11089_),
    .A2(_11244_),
    .B1(_11245_),
    .B2(_11130_),
    .Y(_11246_));
 sky130_fd_sc_hd__a22o_1 _16741_ (.A1(net68),
    .A2(net3546),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[15] ),
    .X(_11247_));
 sky130_fd_sc_hd__a221o_4 _16742_ (.A1(\cs_registers_i.mscratch_q[15] ),
    .A2(net3540),
    .B1(_11063_),
    .B2(\cs_registers_i.dcsr_q[15] ),
    .C1(_11247_),
    .X(_11248_));
 sky130_fd_sc_hd__a21oi_1 _16743_ (.A1(\cs_registers_i.mtval_q[15] ),
    .A2(net3539),
    .B1(_11052_),
    .Y(_11249_));
 sky130_fd_sc_hd__a22oi_2 _16744_ (.A1(\cs_registers_i.csr_mtvec_o[15] ),
    .A2(net3550),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .Y(_11250_));
 sky130_fd_sc_hd__a22oi_1 _16745_ (.A1(\cs_registers_i.dscratch0_q[15] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[15] ),
    .Y(_11251_));
 sky130_fd_sc_hd__nand3_2 _16746_ (.A(_11249_),
    .B(_11250_),
    .C(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__a211oi_4 _16747_ (.A1(_10993_),
    .A2(_11246_),
    .B1(_11248_),
    .C1(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__nor3_1 _16748_ (.A(net3590),
    .B(_10991_),
    .C(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__a21oi_4 _16749_ (.A1(net3590),
    .A2(_10965_),
    .B1(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_818 ();
 sky130_fd_sc_hd__nand2_1 _16751_ (.A(_11118_),
    .B(_11238_),
    .Y(_11257_));
 sky130_fd_sc_hd__a21oi_1 _16752_ (.A1(_11240_),
    .A2(_11257_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .Y(_11258_));
 sky130_fd_sc_hd__a221oi_1 _16753_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_11239_),
    .B1(_11255_),
    .B2(_11120_),
    .C1(_11258_),
    .Y(_00023_));
 sky130_fd_sc_hd__a221o_4 _16754_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(_11098_),
    .B1(_11057_),
    .B2(\cs_registers_i.dscratch0_q[16] ),
    .C1(_11052_),
    .X(_11259_));
 sky130_fd_sc_hd__a22oi_1 _16755_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1872] ),
    .Y(_11260_));
 sky130_fd_sc_hd__a22oi_2 _16756_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1904] ),
    .Y(_11261_));
 sky130_fd_sc_hd__o22ai_4 _16757_ (.A1(_11130_),
    .A2(_11260_),
    .B1(_11261_),
    .B2(_11089_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand2_4 _16758_ (.A(_10993_),
    .B(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__a222oi_1 _16759_ (.A1(net130),
    .A2(_11104_),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[16] ),
    .C1(net69),
    .C2(_11070_),
    .Y(_11264_));
 sky130_fd_sc_hd__a22oi_2 _16760_ (.A1(\cs_registers_i.mtval_q[16] ),
    .A2(net3539),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .Y(_11265_));
 sky130_fd_sc_hd__a22oi_2 _16761_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(net3550),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[16] ),
    .Y(_11266_));
 sky130_fd_sc_hd__nand4_1 _16762_ (.A(_11263_),
    .B(_11264_),
    .C(_11265_),
    .D(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__a211oi_4 _16763_ (.A1(\cs_registers_i.dscratch1_q[16] ),
    .A2(_11059_),
    .B1(_11259_),
    .C1(_11267_),
    .Y(_11268_));
 sky130_fd_sc_hd__nor3_1 _16764_ (.A(net3588),
    .B(_10991_),
    .C(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__a21oi_4 _16765_ (.A1(net3588),
    .A2(_10965_),
    .B1(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_817 ();
 sky130_fd_sc_hd__nand4_1 _16767_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .D(_11237_),
    .Y(_11272_));
 sky130_fd_sc_hd__nor2_1 _16768_ (.A(_11112_),
    .B(_11272_),
    .Y(_11273_));
 sky130_fd_sc_hd__a211oi_1 _16769_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_11239_),
    .B1(_11115_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .Y(_11274_));
 sky130_fd_sc_hd__a211oi_1 _16770_ (.A1(_11120_),
    .A2(_11270_),
    .B1(_11273_),
    .C1(_11274_),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_1 _16771_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .Y(_11275_));
 sky130_fd_sc_hd__nor2_1 _16772_ (.A(_11275_),
    .B(_11272_),
    .Y(_11276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_813 ();
 sky130_fd_sc_hd__a22oi_2 _16777_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1873] ),
    .Y(_11281_));
 sky130_fd_sc_hd__a22oi_2 _16778_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1905] ),
    .Y(_11282_));
 sky130_fd_sc_hd__o22ai_4 _16779_ (.A1(_11130_),
    .A2(_11281_),
    .B1(_11282_),
    .B2(_11089_),
    .Y(_11283_));
 sky130_fd_sc_hd__a22oi_2 _16780_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(net3550),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[17] ),
    .Y(_11284_));
 sky130_fd_sc_hd__a22oi_1 _16781_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(_11098_),
    .B1(_11076_),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .Y(_11285_));
 sky130_fd_sc_hd__a22oi_1 _16782_ (.A1(net136),
    .A2(_11104_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[17] ),
    .Y(_11286_));
 sky130_fd_sc_hd__a22oi_1 _16783_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(net3540),
    .B1(_10595_),
    .B2(\cs_registers_i.mstatus_q[1] ),
    .Y(_11287_));
 sky130_fd_sc_hd__nand4_1 _16784_ (.A(_11284_),
    .B(_11285_),
    .C(_11286_),
    .D(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__nand2_1 _16785_ (.A(\cs_registers_i.dscratch1_q[17] ),
    .B(_11059_),
    .Y(_11289_));
 sky130_fd_sc_hd__a221oi_1 _16786_ (.A1(net70),
    .A2(_11070_),
    .B1(_11057_),
    .B2(\cs_registers_i.dscratch0_q[17] ),
    .C1(_11052_),
    .Y(_11290_));
 sky130_fd_sc_hd__nand2_2 _16787_ (.A(_11289_),
    .B(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__a211oi_4 _16788_ (.A1(_10993_),
    .A2(_11283_),
    .B1(_11288_),
    .C1(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__nor3_1 _16789_ (.A(net3613),
    .B(_10991_),
    .C(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__a21oi_4 _16790_ (.A1(net3613),
    .A2(_10965_),
    .B1(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_812 ();
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(_11118_),
    .B(_11272_),
    .Y(_11296_));
 sky130_fd_sc_hd__a21oi_1 _16793_ (.A1(_11240_),
    .A2(_11296_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .Y(_11297_));
 sky130_fd_sc_hd__a221oi_1 _16794_ (.A1(_11118_),
    .A2(_11276_),
    .B1(_11294_),
    .B2(_11120_),
    .C1(_11297_),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_1 _16795_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .Y(_11298_));
 sky130_fd_sc_hd__o21ai_0 _16796_ (.A1(_11112_),
    .A2(_11276_),
    .B1(_11240_),
    .Y(_11299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_811 ();
 sky130_fd_sc_hd__nand2_1 _16798_ (.A(\cs_registers_i.mhpmcounter[1874] ),
    .B(_10610_),
    .Y(_11301_));
 sky130_fd_sc_hd__o21ai_2 _16799_ (.A1(_11298_),
    .A2(_10996_),
    .B1(_11301_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand2_8 _16800_ (.A(_11001_),
    .B(_10580_),
    .Y(_11303_));
 sky130_fd_sc_hd__a22oi_1 _16801_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1906] ),
    .Y(_11304_));
 sky130_fd_sc_hd__nor2_1 _16802_ (.A(_11303_),
    .B(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__a21oi_4 _16803_ (.A1(_11002_),
    .A2(_11302_),
    .B1(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__nor2_4 _16804_ (.A(_11036_),
    .B(_10602_),
    .Y(_11307_));
 sky130_fd_sc_hd__a221oi_1 _16805_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(_11307_),
    .B1(_11024_),
    .B2(\cs_registers_i.dscratch0_q[18] ),
    .C1(_11015_),
    .Y(_11308_));
 sky130_fd_sc_hd__nor4_1 _16806_ (.A(_10576_),
    .B(_10556_),
    .C(_10560_),
    .D(_11018_),
    .Y(_11309_));
 sky130_fd_sc_hd__a22o_1 _16807_ (.A1(\cs_registers_i.csr_mepc_o[18] ),
    .A2(_11035_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[18] ),
    .X(_11310_));
 sky130_fd_sc_hd__a221oi_4 _16808_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_11029_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .C1(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__nor2_4 _16809_ (.A(_11026_),
    .B(_10602_),
    .Y(_11312_));
 sky130_fd_sc_hd__a222oi_1 _16810_ (.A1(\cs_registers_i.mscratch_q[18] ),
    .A2(_11028_),
    .B1(_11032_),
    .B2(net71),
    .C1(_11312_),
    .C2(net137),
    .Y(_11313_));
 sky130_fd_sc_hd__o2111ai_2 _16811_ (.A1(_11093_),
    .A2(_11306_),
    .B1(_11308_),
    .C1(_11311_),
    .D1(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__a21oi_4 _16812_ (.A1(\cs_registers_i.dscratch1_q[18] ),
    .A2(_11023_),
    .B1(_11314_),
    .Y(_11315_));
 sky130_fd_sc_hd__nor2_1 _16813_ (.A(_10991_),
    .B(_11315_),
    .Y(_11316_));
 sky130_fd_sc_hd__nor2_4 _16814_ (.A(_08008_),
    .B(_10991_),
    .Y(_11317_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(_09663_),
    .B(_11317_),
    .Y(_11318_));
 sky130_fd_sc_hd__o21ai_4 _16816_ (.A1(_09663_),
    .A2(_11316_),
    .B1(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_810 ();
 sky130_fd_sc_hd__a32o_1 _16818_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .A2(_11118_),
    .A3(_11276_),
    .B1(_11319_),
    .B2(_11120_),
    .X(_11321_));
 sky130_fd_sc_hd__a21oi_1 _16819_ (.A1(_11298_),
    .A2(_11299_),
    .B1(_11321_),
    .Y(_00026_));
 sky130_fd_sc_hd__a22o_4 _16820_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1875] ),
    .X(_11322_));
 sky130_fd_sc_hd__a22o_1 _16821_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1907] ),
    .X(_11323_));
 sky130_fd_sc_hd__a22oi_2 _16822_ (.A1(_11002_),
    .A2(_11322_),
    .B1(_11323_),
    .B2(_11004_),
    .Y(_11324_));
 sky130_fd_sc_hd__a221oi_1 _16823_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(_11307_),
    .B1(_11024_),
    .B2(\cs_registers_i.dscratch0_q[19] ),
    .C1(_11015_),
    .Y(_11325_));
 sky130_fd_sc_hd__a22o_1 _16824_ (.A1(\cs_registers_i.csr_mepc_o[19] ),
    .A2(_11035_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[19] ),
    .X(_11326_));
 sky130_fd_sc_hd__a221oi_2 _16825_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_11029_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[19] ),
    .C1(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__a222oi_1 _16826_ (.A1(\cs_registers_i.mscratch_q[19] ),
    .A2(_11028_),
    .B1(_11032_),
    .B2(net72),
    .C1(_11312_),
    .C2(net138),
    .Y(_11328_));
 sky130_fd_sc_hd__o2111ai_2 _16827_ (.A1(_11093_),
    .A2(_11324_),
    .B1(_11325_),
    .C1(_11327_),
    .D1(_11328_),
    .Y(_11329_));
 sky130_fd_sc_hd__a21oi_4 _16828_ (.A1(\cs_registers_i.dscratch1_q[19] ),
    .A2(_11023_),
    .B1(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__nor2_1 _16829_ (.A(_10991_),
    .B(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__nand2_1 _16830_ (.A(_09593_),
    .B(_11317_),
    .Y(_11332_));
 sky130_fd_sc_hd__o21ai_4 _16831_ (.A1(_09593_),
    .A2(_11331_),
    .B1(_11332_),
    .Y(_11333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_809 ();
 sky130_fd_sc_hd__and3_4 _16833_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .X(_11335_));
 sky130_fd_sc_hd__nand3_1 _16834_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .C(_11335_),
    .Y(_11336_));
 sky130_fd_sc_hd__nor2_1 _16835_ (.A(_11241_),
    .B(_11336_),
    .Y(_11337_));
 sky130_fd_sc_hd__and3_1 _16836_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .B(_11113_),
    .C(_11337_),
    .X(_11338_));
 sky130_fd_sc_hd__a211oi_1 _16837_ (.A1(_11113_),
    .A2(_11337_),
    .B1(_11115_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .Y(_11339_));
 sky130_fd_sc_hd__a211oi_1 _16838_ (.A1(_11115_),
    .A2(_11333_),
    .B1(_11338_),
    .C1(_11339_),
    .Y(_00027_));
 sky130_fd_sc_hd__nand2b_1 _16839_ (.A_N(\cs_registers_i.mcountinhibit_q[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .Y(_11340_));
 sky130_fd_sc_hd__a21oi_1 _16840_ (.A1(_11087_),
    .A2(_11340_),
    .B1(_11091_),
    .Y(_11341_));
 sky130_fd_sc_hd__nor2_4 _16841_ (.A(_10585_),
    .B(_10565_),
    .Y(_11342_));
 sky130_fd_sc_hd__a222oi_1 _16842_ (.A1(\cs_registers_i.mcause_q[1] ),
    .A2(_10613_),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .C1(_11342_),
    .C2(\cs_registers_i.dcsr_q[1] ),
    .Y(_11343_));
 sky130_fd_sc_hd__a22oi_1 _16843_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1857] ),
    .Y(_11344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_808 ();
 sky130_fd_sc_hd__a22oi_2 _16845_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1889] ),
    .Y(_11346_));
 sky130_fd_sc_hd__o22ai_2 _16846_ (.A1(_11130_),
    .A2(_11344_),
    .B1(_11346_),
    .B2(_11089_),
    .Y(_11347_));
 sky130_fd_sc_hd__nand2_4 _16847_ (.A(_11085_),
    .B(_11347_),
    .Y(_11348_));
 sky130_fd_sc_hd__a22o_1 _16848_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(net3539),
    .B1(net3552),
    .B2(net73),
    .X(_11349_));
 sky130_fd_sc_hd__a221oi_4 _16849_ (.A1(\cs_registers_i.mscratch_q[1] ),
    .A2(net3540),
    .B1(_11221_),
    .B2(\cs_registers_i.csr_depc_o[1] ),
    .C1(_11349_),
    .Y(_11350_));
 sky130_fd_sc_hd__a22oi_1 _16850_ (.A1(\cs_registers_i.dscratch1_q[1] ),
    .A2(_11227_),
    .B1(_11228_),
    .B2(\cs_registers_i.dscratch0_q[1] ),
    .Y(_11351_));
 sky130_fd_sc_hd__and4_4 _16851_ (.A(_11343_),
    .B(_11348_),
    .C(_11350_),
    .D(_11351_),
    .X(_11352_));
 sky130_fd_sc_hd__nor3_1 _16852_ (.A(net3597),
    .B(_10991_),
    .C(_11352_),
    .Y(_11353_));
 sky130_fd_sc_hd__a21oi_4 _16853_ (.A1(net3597),
    .A2(_10965_),
    .B1(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_807 ();
 sky130_fd_sc_hd__a32oi_1 _16855_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A3(_11113_),
    .B1(_11120_),
    .B2(_11354_),
    .Y(_11356_));
 sky130_fd_sc_hd__o21a_1 _16856_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A2(_11341_),
    .B1(_11356_),
    .X(_00028_));
 sky130_fd_sc_hd__a22o_4 _16857_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1876] ),
    .X(_11357_));
 sky130_fd_sc_hd__a22o_1 _16858_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1908] ),
    .X(_11358_));
 sky130_fd_sc_hd__a22oi_2 _16859_ (.A1(_11002_),
    .A2(_11357_),
    .B1(_11358_),
    .B2(_11004_),
    .Y(_11359_));
 sky130_fd_sc_hd__a22o_1 _16860_ (.A1(\cs_registers_i.mscratch_q[20] ),
    .A2(_11028_),
    .B1(_11312_),
    .B2(net139),
    .X(_11360_));
 sky130_fd_sc_hd__a221oi_2 _16861_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_11029_),
    .B1(_11035_),
    .B2(\cs_registers_i.csr_mepc_o[20] ),
    .C1(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__a22o_1 _16862_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(_11307_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[20] ),
    .X(_11362_));
 sky130_fd_sc_hd__a221oi_2 _16863_ (.A1(net74),
    .A2(_11032_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .C1(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__o21bai_4 _16864_ (.A1(_10576_),
    .A2(_11036_),
    .B1_N(_11015_),
    .Y(_11364_));
 sky130_fd_sc_hd__a221oi_2 _16865_ (.A1(\cs_registers_i.dscratch1_q[20] ),
    .A2(_11023_),
    .B1(_11024_),
    .B2(\cs_registers_i.dscratch0_q[20] ),
    .C1(_11364_),
    .Y(_11365_));
 sky130_fd_sc_hd__o2111ai_4 _16866_ (.A1(_11093_),
    .A2(_11359_),
    .B1(_11361_),
    .C1(_11363_),
    .D1(_11365_),
    .Y(_11366_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(_10964_),
    .B(_11366_),
    .Y(_11367_));
 sky130_fd_sc_hd__nand2_2 _16868_ (.A(_09797_),
    .B(_11367_),
    .Y(_11368_));
 sky130_fd_sc_hd__o21ai_4 _16869_ (.A1(_09797_),
    .A2(_10965_),
    .B1(_11368_),
    .Y(_11369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_806 ();
 sky130_fd_sc_hd__nand4_1 _16871_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .C(_11217_),
    .D(_11335_),
    .Y(_11371_));
 sky130_fd_sc_hd__nand3_1 _16872_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .C(_11157_),
    .Y(_11372_));
 sky130_fd_sc_hd__nor2_1 _16873_ (.A(_11371_),
    .B(_11372_),
    .Y(_11373_));
 sky130_fd_sc_hd__and3_4 _16874_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .B(_11113_),
    .C(_11373_),
    .X(_11374_));
 sky130_fd_sc_hd__o31ai_1 _16875_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11371_),
    .A3(_11372_),
    .B1(_11118_),
    .Y(_11375_));
 sky130_fd_sc_hd__a21oi_1 _16876_ (.A1(_11240_),
    .A2(_11375_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .Y(_11376_));
 sky130_fd_sc_hd__a211oi_1 _16877_ (.A1(_11120_),
    .A2(_11369_),
    .B1(_11374_),
    .C1(_11376_),
    .Y(_00029_));
 sky130_fd_sc_hd__a22oi_1 _16878_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1877] ),
    .Y(_11377_));
 sky130_fd_sc_hd__a22oi_2 _16879_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1909] ),
    .Y(_11378_));
 sky130_fd_sc_hd__o22ai_4 _16880_ (.A1(_11130_),
    .A2(_11377_),
    .B1(_11378_),
    .B2(_11089_),
    .Y(_11379_));
 sky130_fd_sc_hd__a22oi_2 _16881_ (.A1(\cs_registers_i.csr_mtvec_o[21] ),
    .A2(net3550),
    .B1(_10625_),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .Y(_11380_));
 sky130_fd_sc_hd__a22oi_1 _16882_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(_11098_),
    .B1(_11076_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .Y(_11381_));
 sky130_fd_sc_hd__a22oi_2 _16883_ (.A1(net140),
    .A2(_11104_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[21] ),
    .Y(_11382_));
 sky130_fd_sc_hd__a22oi_1 _16884_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(net3540),
    .B1(_10595_),
    .B2(\cs_registers_i.csr_mstatus_tw_o ),
    .Y(_11383_));
 sky130_fd_sc_hd__nand4_1 _16885_ (.A(_11380_),
    .B(_11381_),
    .C(_11382_),
    .D(_11383_),
    .Y(_11384_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(\cs_registers_i.dscratch1_q[21] ),
    .B(_11059_),
    .Y(_11385_));
 sky130_fd_sc_hd__a221oi_1 _16887_ (.A1(net75),
    .A2(_11070_),
    .B1(_11057_),
    .B2(\cs_registers_i.dscratch0_q[21] ),
    .C1(_11052_),
    .Y(_11386_));
 sky130_fd_sc_hd__nand2_2 _16888_ (.A(_11385_),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__a211oi_4 _16889_ (.A1(_10993_),
    .A2(_11379_),
    .B1(_11384_),
    .C1(_11387_),
    .Y(_11388_));
 sky130_fd_sc_hd__nor3_1 _16890_ (.A(_09730_),
    .B(_10991_),
    .C(_11388_),
    .Y(_11389_));
 sky130_fd_sc_hd__a21oi_4 _16891_ (.A1(_09730_),
    .A2(_10965_),
    .B1(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_805 ();
 sky130_fd_sc_hd__nor3_1 _16893_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .B(_11115_),
    .C(_11374_),
    .Y(_11392_));
 sky130_fd_sc_hd__a21o_1 _16894_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(_11374_),
    .B1(_11392_),
    .X(_11393_));
 sky130_fd_sc_hd__a21oi_1 _16895_ (.A1(_11120_),
    .A2(net3494),
    .B1(_11393_),
    .Y(_00030_));
 sky130_fd_sc_hd__a22o_1 _16896_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1878] ),
    .X(_11394_));
 sky130_fd_sc_hd__inv_1 _16897_ (.A(\cs_registers_i.mhpmcounter[1910] ),
    .Y(_11395_));
 sky130_fd_sc_hd__nand2_1 _16898_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .B(net3581),
    .Y(_11396_));
 sky130_fd_sc_hd__o21ai_0 _16899_ (.A1(_11395_),
    .A2(_11009_),
    .B1(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__a22oi_2 _16900_ (.A1(_11002_),
    .A2(_11394_),
    .B1(_11397_),
    .B2(_11004_),
    .Y(_11398_));
 sky130_fd_sc_hd__a221oi_1 _16901_ (.A1(net76),
    .A2(_11032_),
    .B1(_11023_),
    .B2(\cs_registers_i.dscratch1_q[22] ),
    .C1(_11015_),
    .Y(_11399_));
 sky130_fd_sc_hd__a22o_1 _16902_ (.A1(\cs_registers_i.mscratch_q[22] ),
    .A2(_11028_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[22] ),
    .X(_11400_));
 sky130_fd_sc_hd__a221oi_4 _16903_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_11029_),
    .B1(_11035_),
    .B2(\cs_registers_i.csr_mepc_o[22] ),
    .C1(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__a222oi_1 _16904_ (.A1(net141),
    .A2(_11312_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .C1(_11307_),
    .C2(\cs_registers_i.mie_q[6] ),
    .Y(_11402_));
 sky130_fd_sc_hd__o2111ai_2 _16905_ (.A1(_11093_),
    .A2(_11398_),
    .B1(_11399_),
    .C1(_11401_),
    .D1(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__a21oi_4 _16906_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_11024_),
    .B1(_11403_),
    .Y(_11404_));
 sky130_fd_sc_hd__o21ai_2 _16907_ (.A1(_10991_),
    .A2(_11404_),
    .B1(net437),
    .Y(_11405_));
 sky130_fd_sc_hd__o21ai_4 _16908_ (.A1(net437),
    .A2(_10965_),
    .B1(_11405_),
    .Y(_11406_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_804 ();
 sky130_fd_sc_hd__a211oi_1 _16910_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(_11374_),
    .B1(_11120_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .Y(_11408_));
 sky130_fd_sc_hd__a31o_1 _16911_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A3(_11374_),
    .B1(_11408_),
    .X(_11409_));
 sky130_fd_sc_hd__a21oi_1 _16912_ (.A1(_11115_),
    .A2(net3493),
    .B1(_11409_),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _16913_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .Y(_11410_));
 sky130_fd_sc_hd__nand4_1 _16914_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .D(_11373_),
    .Y(_11411_));
 sky130_fd_sc_hd__nor2_1 _16915_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__o21ai_0 _16916_ (.A1(_11112_),
    .A2(_11412_),
    .B1(_11240_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(\cs_registers_i.mhpmcounter[1879] ),
    .B(_10610_),
    .Y(_11414_));
 sky130_fd_sc_hd__o21ai_2 _16918_ (.A1(_11410_),
    .A2(_10996_),
    .B1(_11414_),
    .Y(_11415_));
 sky130_fd_sc_hd__a22o_1 _16919_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1911] ),
    .X(_11416_));
 sky130_fd_sc_hd__a22oi_2 _16920_ (.A1(_11002_),
    .A2(_11415_),
    .B1(_11416_),
    .B2(_11004_),
    .Y(_11417_));
 sky130_fd_sc_hd__a221oi_1 _16921_ (.A1(net77),
    .A2(_11032_),
    .B1(_11023_),
    .B2(\cs_registers_i.dscratch1_q[23] ),
    .C1(_11015_),
    .Y(_11418_));
 sky130_fd_sc_hd__a22o_1 _16922_ (.A1(\cs_registers_i.mscratch_q[23] ),
    .A2(_11028_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .X(_11419_));
 sky130_fd_sc_hd__a221oi_4 _16923_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_11029_),
    .B1(_11035_),
    .B2(\cs_registers_i.csr_mepc_o[23] ),
    .C1(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__a222oi_1 _16924_ (.A1(net142),
    .A2(_11312_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C1(_11307_),
    .C2(\cs_registers_i.mie_q[7] ),
    .Y(_11421_));
 sky130_fd_sc_hd__o2111ai_2 _16925_ (.A1(_11093_),
    .A2(_11417_),
    .B1(_11418_),
    .C1(_11420_),
    .D1(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__a21oi_4 _16926_ (.A1(\cs_registers_i.dscratch0_q[23] ),
    .A2(_11024_),
    .B1(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__nor2_1 _16927_ (.A(_10991_),
    .B(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(_09907_),
    .B(_11317_),
    .Y(_11425_));
 sky130_fd_sc_hd__o21ai_4 _16929_ (.A1(_09907_),
    .A2(_11424_),
    .B1(_11425_),
    .Y(_11426_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_803 ();
 sky130_fd_sc_hd__and3_4 _16931_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .B(_11118_),
    .C(_11412_),
    .X(_11428_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_11120_),
    .A2(net3492),
    .B1(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__a21oi_1 _16933_ (.A1(_11410_),
    .A2(_11413_),
    .B1(_11429_),
    .Y(_00032_));
 sky130_fd_sc_hd__a221o_4 _16934_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(_11098_),
    .B1(net3548),
    .B2(\cs_registers_i.dscratch0_q[24] ),
    .C1(_11052_),
    .X(_11430_));
 sky130_fd_sc_hd__a22oi_2 _16935_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1880] ),
    .Y(_11431_));
 sky130_fd_sc_hd__a22oi_2 _16936_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1912] ),
    .Y(_11432_));
 sky130_fd_sc_hd__o22ai_4 _16937_ (.A1(_11130_),
    .A2(_11431_),
    .B1(_11432_),
    .B2(_11089_),
    .Y(_11433_));
 sky130_fd_sc_hd__nand2_2 _16938_ (.A(_10993_),
    .B(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__a222oi_1 _16939_ (.A1(net143),
    .A2(_11104_),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[24] ),
    .C1(net78),
    .C2(_11070_),
    .Y(_11435_));
 sky130_fd_sc_hd__a22oi_2 _16940_ (.A1(\cs_registers_i.mtval_q[24] ),
    .A2(net3539),
    .B1(_11076_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .Y(_11436_));
 sky130_fd_sc_hd__a22oi_2 _16941_ (.A1(\cs_registers_i.csr_mtvec_o[24] ),
    .A2(net3550),
    .B1(_10625_),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .Y(_11437_));
 sky130_fd_sc_hd__nand4_1 _16942_ (.A(_11434_),
    .B(_11435_),
    .C(_11436_),
    .D(_11437_),
    .Y(_11438_));
 sky130_fd_sc_hd__a211oi_4 _16943_ (.A1(\cs_registers_i.dscratch1_q[24] ),
    .A2(net3547),
    .B1(_11430_),
    .C1(_11438_),
    .Y(_11439_));
 sky130_fd_sc_hd__nor3_1 _16944_ (.A(_09986_),
    .B(_10991_),
    .C(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__a21oi_4 _16945_ (.A1(_09986_),
    .A2(_10965_),
    .B1(_11440_),
    .Y(_11441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_802 ();
 sky130_fd_sc_hd__nor3_1 _16947_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .B(_11120_),
    .C(_11428_),
    .Y(_11443_));
 sky130_fd_sc_hd__and2_4 _16948_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .B(_11428_),
    .X(_11444_));
 sky130_fd_sc_hd__a211oi_1 _16949_ (.A1(_11115_),
    .A2(net3483),
    .B1(_11443_),
    .C1(_11444_),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_2 _16950_ (.A(\cs_registers_i.mhpmcounter[1881] ),
    .Y(_11445_));
 sky130_fd_sc_hd__nand2_1 _16951_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .B(net3581),
    .Y(_11446_));
 sky130_fd_sc_hd__o21ai_2 _16952_ (.A1(_11445_),
    .A2(_11009_),
    .B1(_11446_),
    .Y(_11447_));
 sky130_fd_sc_hd__a22o_1 _16953_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1913] ),
    .X(_11448_));
 sky130_fd_sc_hd__a22oi_2 _16954_ (.A1(_11002_),
    .A2(_11447_),
    .B1(_11448_),
    .B2(_11004_),
    .Y(_11449_));
 sky130_fd_sc_hd__a221oi_1 _16955_ (.A1(net79),
    .A2(_11032_),
    .B1(_11023_),
    .B2(\cs_registers_i.dscratch1_q[25] ),
    .C1(_11015_),
    .Y(_11450_));
 sky130_fd_sc_hd__a22o_1 _16956_ (.A1(\cs_registers_i.mscratch_q[25] ),
    .A2(_11028_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[25] ),
    .X(_11451_));
 sky130_fd_sc_hd__a221oi_4 _16957_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_11029_),
    .B1(_11035_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .C1(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__a222oi_1 _16958_ (.A1(net144),
    .A2(_11312_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .C1(_11307_),
    .C2(\cs_registers_i.mie_q[9] ),
    .Y(_11453_));
 sky130_fd_sc_hd__o2111ai_2 _16959_ (.A1(_11093_),
    .A2(_11449_),
    .B1(_11450_),
    .C1(_11452_),
    .D1(_11453_),
    .Y(_11454_));
 sky130_fd_sc_hd__a21oi_4 _16960_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(_11024_),
    .B1(_11454_),
    .Y(_11455_));
 sky130_fd_sc_hd__o21ai_1 _16961_ (.A1(_10991_),
    .A2(_11455_),
    .B1(_10098_),
    .Y(_11456_));
 sky130_fd_sc_hd__o21ai_4 _16962_ (.A1(_10098_),
    .A2(_10965_),
    .B1(_11456_),
    .Y(_11457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_801 ();
 sky130_fd_sc_hd__nor3_1 _16964_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .B(_11120_),
    .C(_11444_),
    .Y(_11459_));
 sky130_fd_sc_hd__a21o_1 _16965_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A2(_11444_),
    .B1(_11459_),
    .X(_11460_));
 sky130_fd_sc_hd__a21oi_1 _16966_ (.A1(_11115_),
    .A2(_11457_),
    .B1(_11460_),
    .Y(_00034_));
 sky130_fd_sc_hd__a21oi_1 _16967_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A2(_11444_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .Y(_11461_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(_11202_),
    .B(_11461_),
    .Y(_11462_));
 sky130_fd_sc_hd__nand3_1 _16969_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .C(_11444_),
    .Y(_11463_));
 sky130_fd_sc_hd__a221o_4 _16970_ (.A1(net80),
    .A2(_11070_),
    .B1(net3547),
    .B2(\cs_registers_i.dscratch1_q[26] ),
    .C1(_11052_),
    .X(_11464_));
 sky130_fd_sc_hd__a22oi_2 _16971_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1882] ),
    .Y(_11465_));
 sky130_fd_sc_hd__a22oi_2 _16972_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1914] ),
    .Y(_11466_));
 sky130_fd_sc_hd__o22ai_4 _16973_ (.A1(_11130_),
    .A2(_11465_),
    .B1(_11466_),
    .B2(_11089_),
    .Y(_11467_));
 sky130_fd_sc_hd__nand2_4 _16974_ (.A(_10993_),
    .B(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__a22oi_1 _16975_ (.A1(\cs_registers_i.csr_mepc_o[26] ),
    .A2(_10625_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[26] ),
    .Y(_11469_));
 sky130_fd_sc_hd__a22oi_1 _16976_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[26] ),
    .Y(_11470_));
 sky130_fd_sc_hd__a222oi_1 _16977_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(_11098_),
    .B1(_11104_),
    .B2(net131),
    .C1(_11076_),
    .C2(\cs_registers_i.csr_depc_o[26] ),
    .Y(_11471_));
 sky130_fd_sc_hd__nand4_1 _16978_ (.A(_11468_),
    .B(_11469_),
    .C(_11470_),
    .D(_11471_),
    .Y(_11472_));
 sky130_fd_sc_hd__a211oi_4 _16979_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(net3548),
    .B1(_11464_),
    .C1(_11472_),
    .Y(_11473_));
 sky130_fd_sc_hd__nor2_2 _16980_ (.A(_10991_),
    .B(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__nor2_1 _16981_ (.A(_10173_),
    .B(_11317_),
    .Y(_11475_));
 sky130_fd_sc_hd__a21oi_4 _16982_ (.A1(_10173_),
    .A2(_11474_),
    .B1(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_800 ();
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(_11115_),
    .B(net3482),
    .Y(_11478_));
 sky130_fd_sc_hd__and3_1 _16985_ (.A(_11462_),
    .B(_11463_),
    .C(_11478_),
    .X(_00035_));
 sky130_fd_sc_hd__a221o_4 _16986_ (.A1(net81),
    .A2(_11070_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[27] ),
    .C1(_11052_),
    .X(_11479_));
 sky130_fd_sc_hd__a22oi_2 _16987_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1883] ),
    .Y(_11480_));
 sky130_fd_sc_hd__a22oi_2 _16988_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1915] ),
    .Y(_11481_));
 sky130_fd_sc_hd__o22ai_4 _16989_ (.A1(_11130_),
    .A2(_11480_),
    .B1(_11481_),
    .B2(_11089_),
    .Y(_11482_));
 sky130_fd_sc_hd__nand2_4 _16990_ (.A(_10993_),
    .B(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__a22oi_1 _16991_ (.A1(\cs_registers_i.csr_mepc_o[27] ),
    .A2(_10625_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[27] ),
    .Y(_11484_));
 sky130_fd_sc_hd__a22oi_1 _16992_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[27] ),
    .Y(_11485_));
 sky130_fd_sc_hd__a222oi_1 _16993_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(_11098_),
    .B1(_11104_),
    .B2(net132),
    .C1(_11076_),
    .C2(\cs_registers_i.csr_depc_o[27] ),
    .Y(_11486_));
 sky130_fd_sc_hd__nand4_1 _16994_ (.A(_11483_),
    .B(_11484_),
    .C(_11485_),
    .D(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__a211oi_4 _16995_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_11057_),
    .B1(_11479_),
    .C1(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__nor3_1 _16996_ (.A(_10203_),
    .B(_10991_),
    .C(_11488_),
    .Y(_11489_));
 sky130_fd_sc_hd__a21oi_4 _16997_ (.A1(_10203_),
    .A2(_10965_),
    .B1(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_799 ();
 sky130_fd_sc_hd__nor2_1 _16999_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .B(_11120_),
    .Y(_11492_));
 sky130_fd_sc_hd__mux2_1 _17000_ (.A0(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A1(_11492_),
    .S(_11463_),
    .X(_11493_));
 sky130_fd_sc_hd__a21oi_1 _17001_ (.A1(_11120_),
    .A2(net3481),
    .B1(_11493_),
    .Y(_00036_));
 sky130_fd_sc_hd__a221o_4 _17002_ (.A1(net82),
    .A2(_11070_),
    .B1(net3547),
    .B2(\cs_registers_i.dscratch1_q[28] ),
    .C1(_11052_),
    .X(_11494_));
 sky130_fd_sc_hd__a22oi_2 _17003_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1884] ),
    .Y(_11495_));
 sky130_fd_sc_hd__a22oi_2 _17004_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1916] ),
    .Y(_11496_));
 sky130_fd_sc_hd__o22ai_4 _17005_ (.A1(_11130_),
    .A2(_11495_),
    .B1(_11496_),
    .B2(_11089_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_8 _17006_ (.A(_10993_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__a22oi_1 _17007_ (.A1(\cs_registers_i.csr_mepc_o[28] ),
    .A2(_10625_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[28] ),
    .Y(_11499_));
 sky130_fd_sc_hd__a22oi_1 _17008_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[28] ),
    .Y(_11500_));
 sky130_fd_sc_hd__a222oi_1 _17009_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(_11098_),
    .B1(_11104_),
    .B2(net133),
    .C1(_11076_),
    .C2(\cs_registers_i.csr_depc_o[28] ),
    .Y(_11501_));
 sky130_fd_sc_hd__nand4_1 _17010_ (.A(_11498_),
    .B(_11499_),
    .C(_11500_),
    .D(_11501_),
    .Y(_11502_));
 sky130_fd_sc_hd__a211oi_4 _17011_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(net3548),
    .B1(_11494_),
    .C1(_11502_),
    .Y(_11503_));
 sky130_fd_sc_hd__nor2_2 _17012_ (.A(_10991_),
    .B(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__nor2_1 _17013_ (.A(_10269_),
    .B(_11317_),
    .Y(_11505_));
 sky130_fd_sc_hd__a21oi_4 _17014_ (.A1(_10269_),
    .A2(_11504_),
    .B1(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_798 ();
 sky130_fd_sc_hd__nand4_1 _17016_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .D(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .Y(_11508_));
 sky130_fd_sc_hd__nor3_2 _17017_ (.A(_11410_),
    .B(_11411_),
    .C(_11508_),
    .Y(_11509_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .B(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__nor3_1 _17019_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(net3484),
    .C(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__nand2b_1 _17020_ (.A_N(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11509_),
    .Y(_11512_));
 sky130_fd_sc_hd__a21oi_1 _17021_ (.A1(_11118_),
    .A2(_11512_),
    .B1(_11091_),
    .Y(_11513_));
 sky130_fd_sc_hd__nor2_1 _17022_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .B(_11513_),
    .Y(_11514_));
 sky130_fd_sc_hd__a211oi_1 _17023_ (.A1(_11120_),
    .A2(net3480),
    .B1(_11511_),
    .C1(_11514_),
    .Y(_00037_));
 sky130_fd_sc_hd__o21ai_0 _17024_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11510_),
    .B1(_11118_),
    .Y(_11515_));
 sky130_fd_sc_hd__a21oi_1 _17025_ (.A1(_11240_),
    .A2(_11515_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .Y(_11516_));
 sky130_fd_sc_hd__nand4_1 _17026_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .C(_11113_),
    .D(_11509_),
    .Y(_11517_));
 sky130_fd_sc_hd__a221o_4 _17027_ (.A1(net83),
    .A2(_11070_),
    .B1(net3547),
    .B2(\cs_registers_i.dscratch1_q[29] ),
    .C1(_11052_),
    .X(_11518_));
 sky130_fd_sc_hd__a22oi_2 _17028_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1885] ),
    .Y(_11519_));
 sky130_fd_sc_hd__a22oi_2 _17029_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1917] ),
    .Y(_11520_));
 sky130_fd_sc_hd__o22ai_4 _17030_ (.A1(_11130_),
    .A2(_11519_),
    .B1(_11520_),
    .B2(_11089_),
    .Y(_11521_));
 sky130_fd_sc_hd__nand2_8 _17031_ (.A(_10993_),
    .B(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__a22oi_1 _17032_ (.A1(\cs_registers_i.csr_mepc_o[29] ),
    .A2(_10625_),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[29] ),
    .Y(_11523_));
 sky130_fd_sc_hd__a22oi_1 _17033_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[29] ),
    .Y(_11524_));
 sky130_fd_sc_hd__a222oi_1 _17034_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(_11098_),
    .B1(_11104_),
    .B2(net134),
    .C1(_11076_),
    .C2(\cs_registers_i.csr_depc_o[29] ),
    .Y(_11525_));
 sky130_fd_sc_hd__nand4_1 _17035_ (.A(_11522_),
    .B(_11523_),
    .C(_11524_),
    .D(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__a211oi_4 _17036_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(net3548),
    .B1(_11518_),
    .C1(_11526_),
    .Y(_11527_));
 sky130_fd_sc_hd__nor2_2 _17037_ (.A(_10991_),
    .B(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__nor2_1 _17038_ (.A(_10336_),
    .B(_11317_),
    .Y(_11529_));
 sky130_fd_sc_hd__a21oi_4 _17039_ (.A1(_10336_),
    .A2(_11528_),
    .B1(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_797 ();
 sky130_fd_sc_hd__nand2_1 _17041_ (.A(_11120_),
    .B(net3479),
    .Y(_11532_));
 sky130_fd_sc_hd__nand2_1 _17042_ (.A(_11517_),
    .B(_11532_),
    .Y(_11533_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(_11516_),
    .B(_11533_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _17044_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .Y(_11534_));
 sky130_fd_sc_hd__o21ai_0 _17045_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11534_),
    .B1(_11087_),
    .Y(_11535_));
 sky130_fd_sc_hd__a21oi_1 _17046_ (.A1(_11240_),
    .A2(_11535_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .Y(_11536_));
 sky130_fd_sc_hd__a22o_1 _17047_ (.A1(_11082_),
    .A2(_11120_),
    .B1(_11150_),
    .B2(_11113_),
    .X(_11537_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_11536_),
    .B(_11537_),
    .Y(_00039_));
 sky130_fd_sc_hd__a22oi_2 _17049_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1918] ),
    .Y(_11538_));
 sky130_fd_sc_hd__a22o_1 _17050_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1886] ),
    .X(_11539_));
 sky130_fd_sc_hd__nand2_1 _17051_ (.A(_11002_),
    .B(_11539_),
    .Y(_11540_));
 sky130_fd_sc_hd__o21ai_4 _17052_ (.A1(_11303_),
    .A2(_11538_),
    .B1(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__a22oi_2 _17053_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_11023_),
    .B1(_11024_),
    .B2(\cs_registers_i.dscratch0_q[30] ),
    .Y(_11542_));
 sky130_fd_sc_hd__a211oi_1 _17054_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_11035_),
    .B1(_11030_),
    .C1(_11364_),
    .Y(_11543_));
 sky130_fd_sc_hd__a222oi_1 _17055_ (.A1(net135),
    .A2(_11312_),
    .B1(net3565),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .C1(_11307_),
    .C2(\cs_registers_i.mie_q[14] ),
    .Y(_11544_));
 sky130_fd_sc_hd__a22o_1 _17056_ (.A1(net85),
    .A2(_11032_),
    .B1(_11037_),
    .B2(\cs_registers_i.csr_mtvec_o[30] ),
    .X(_11545_));
 sky130_fd_sc_hd__a221oi_1 _17057_ (.A1(\cs_registers_i.mscratch_q[30] ),
    .A2(_11028_),
    .B1(_11029_),
    .B2(\cs_registers_i.mtval_q[30] ),
    .C1(_11545_),
    .Y(_11546_));
 sky130_fd_sc_hd__nand4_1 _17058_ (.A(_11542_),
    .B(_11543_),
    .C(_11544_),
    .D(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__a21oi_4 _17059_ (.A1(_10993_),
    .A2(_11541_),
    .B1(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__o21ai_1 _17060_ (.A1(_10991_),
    .A2(_11548_),
    .B1(_10452_),
    .Y(_11549_));
 sky130_fd_sc_hd__o21ai_4 _17061_ (.A1(_10452_),
    .A2(_10965_),
    .B1(_11549_),
    .Y(_11550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_796 ();
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .B(_11115_),
    .Y(_11552_));
 sky130_fd_sc_hd__mux2_1 _17064_ (.A0(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A1(_11552_),
    .S(_11517_),
    .X(_11553_));
 sky130_fd_sc_hd__a21oi_1 _17065_ (.A1(_11120_),
    .A2(_11550_),
    .B1(_11553_),
    .Y(_00040_));
 sky130_fd_sc_hd__a22oi_2 _17066_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(net3581),
    .B1(net3580),
    .B2(\cs_registers_i.mhpmcounter[1919] ),
    .Y(_11554_));
 sky130_fd_sc_hd__a22oi_2 _17067_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1887] ),
    .Y(_11555_));
 sky130_fd_sc_hd__o22ai_4 _17068_ (.A1(_11089_),
    .A2(_11554_),
    .B1(_11555_),
    .B2(_11130_),
    .Y(_11556_));
 sky130_fd_sc_hd__a22o_1 _17069_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(net3550),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .X(_11557_));
 sky130_fd_sc_hd__a221o_4 _17070_ (.A1(\cs_registers_i.mcause_q[5] ),
    .A2(_10613_),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[31] ),
    .C1(_11557_),
    .X(_11558_));
 sky130_fd_sc_hd__a21oi_1 _17071_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(net3539),
    .B1(_11052_),
    .Y(_11559_));
 sky130_fd_sc_hd__a22oi_1 _17072_ (.A1(net86),
    .A2(_11070_),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[31] ),
    .Y(_11560_));
 sky130_fd_sc_hd__a22oi_2 _17073_ (.A1(\cs_registers_i.dscratch0_q[31] ),
    .A2(net3548),
    .B1(net3547),
    .B2(\cs_registers_i.dscratch1_q[31] ),
    .Y(_11561_));
 sky130_fd_sc_hd__nand3_2 _17074_ (.A(_11559_),
    .B(_11560_),
    .C(_11561_),
    .Y(_11562_));
 sky130_fd_sc_hd__a211oi_4 _17075_ (.A1(_10993_),
    .A2(_11556_),
    .B1(_11558_),
    .C1(_11562_),
    .Y(_11563_));
 sky130_fd_sc_hd__nor3_1 _17076_ (.A(net3587),
    .B(_10991_),
    .C(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__a21oi_4 _17077_ (.A1(net3587),
    .A2(_10965_),
    .B1(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_795 ();
 sky130_fd_sc_hd__and4_4 _17079_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .D(_11509_),
    .X(_11567_));
 sky130_fd_sc_hd__a21o_1 _17080_ (.A1(_11113_),
    .A2(_11567_),
    .B1(_11120_),
    .X(_11568_));
 sky130_fd_sc_hd__nand3_1 _17081_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .B(_11113_),
    .C(_11567_),
    .Y(_11569_));
 sky130_fd_sc_hd__o21ai_0 _17082_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A2(_11568_),
    .B1(_11569_),
    .Y(_11570_));
 sky130_fd_sc_hd__a21oi_1 _17083_ (.A1(_11115_),
    .A2(_11565_),
    .B1(_11570_),
    .Y(_00041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_794 ();
 sky130_fd_sc_hd__nand2_1 _17085_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .B(_11567_),
    .Y(_11572_));
 sky130_fd_sc_hd__nand4_1 _17086_ (.A(net3581),
    .B(_10581_),
    .C(_11085_),
    .D(net3501),
    .Y(_11573_));
 sky130_fd_sc_hd__and2_4 _17087_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(_11573_),
    .X(_11574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_792 ();
 sky130_fd_sc_hd__nor3_1 _17090_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .B(_11572_),
    .C(_11574_),
    .Y(_11577_));
 sky130_fd_sc_hd__a21oi_1 _17091_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A2(_11572_),
    .B1(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__nor3_2 _17092_ (.A(_10996_),
    .B(_11089_),
    .C(_11086_),
    .Y(_11579_));
 sky130_fd_sc_hd__nor2_4 _17093_ (.A(_11113_),
    .B(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_790 ();
 sky130_fd_sc_hd__nor2_1 _17096_ (.A(_11042_),
    .B(net3491),
    .Y(_11583_));
 sky130_fd_sc_hd__a21oi_1 _17097_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A2(_11580_),
    .B1(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__o21ai_0 _17098_ (.A1(_11147_),
    .A2(_11578_),
    .B1(_11584_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand3_2 _17099_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .C(_11567_),
    .Y(_11585_));
 sky130_fd_sc_hd__nor3_1 _17100_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .B(_11574_),
    .C(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__a21oi_1 _17101_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(_11585_),
    .B1(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__nor2_1 _17102_ (.A(_11354_),
    .B(net3491),
    .Y(_11588_));
 sky130_fd_sc_hd__a21oi_1 _17103_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(_11580_),
    .B1(_11588_),
    .Y(_11589_));
 sky130_fd_sc_hd__o21ai_0 _17104_ (.A1(_11147_),
    .A2(_11587_),
    .B1(_11589_),
    .Y(_00043_));
 sky130_fd_sc_hd__and3_4 _17105_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .C(_11567_),
    .X(_11590_));
 sky130_fd_sc_hd__nand2_1 _17106_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .B(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__nor3_1 _17107_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .B(_11574_),
    .C(_11591_),
    .Y(_11592_));
 sky130_fd_sc_hd__a21oi_1 _17108_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(_11591_),
    .B1(_11592_),
    .Y(_11593_));
 sky130_fd_sc_hd__nor2_1 _17109_ (.A(_11082_),
    .B(net3491),
    .Y(_11594_));
 sky130_fd_sc_hd__a21oi_1 _17110_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(_11580_),
    .B1(_11594_),
    .Y(_11595_));
 sky130_fd_sc_hd__o21ai_0 _17111_ (.A1(_11147_),
    .A2(_11593_),
    .B1(_11595_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand3_1 _17112_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .C(_11590_),
    .Y(_11596_));
 sky130_fd_sc_hd__nor3_1 _17113_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .B(_11574_),
    .C(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__a21oi_1 _17114_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(_11596_),
    .B1(_11597_),
    .Y(_11598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_789 ();
 sky130_fd_sc_hd__a22o_1 _17116_ (.A1(\cs_registers_i.mcause_q[3] ),
    .A2(_10613_),
    .B1(_10595_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .X(_11600_));
 sky130_fd_sc_hd__a221oi_4 _17117_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(net3540),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .C1(_11600_),
    .Y(_11601_));
 sky130_fd_sc_hd__a22o_1 _17118_ (.A1(\cs_registers_i.mie_q[17] ),
    .A2(_10620_),
    .B1(_11221_),
    .B2(\cs_registers_i.csr_depc_o[3] ),
    .X(_11602_));
 sky130_fd_sc_hd__a221oi_2 _17119_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(net3539),
    .B1(_10624_),
    .B2(net146),
    .C1(_11602_),
    .Y(_11603_));
 sky130_fd_sc_hd__a22oi_2 _17120_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1891] ),
    .Y(_11604_));
 sky130_fd_sc_hd__a22oi_1 _17121_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1859] ),
    .Y(_11605_));
 sky130_fd_sc_hd__o22ai_2 _17122_ (.A1(_11089_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(_11130_),
    .Y(_11606_));
 sky130_fd_sc_hd__a221o_1 _17123_ (.A1(net87),
    .A2(net3552),
    .B1(_11228_),
    .B2(\cs_registers_i.dscratch0_q[3] ),
    .C1(net3551),
    .X(_11607_));
 sky130_fd_sc_hd__a21oi_1 _17124_ (.A1(_11085_),
    .A2(_11606_),
    .B1(_11607_),
    .Y(_11608_));
 sky130_fd_sc_hd__nand2_1 _17125_ (.A(\cs_registers_i.dscratch1_q[3] ),
    .B(_11227_),
    .Y(_11609_));
 sky130_fd_sc_hd__nand4_1 _17126_ (.A(_11601_),
    .B(_11603_),
    .C(_11608_),
    .D(_11609_),
    .Y(_11610_));
 sky130_fd_sc_hd__nor2_1 _17127_ (.A(net3599),
    .B(_11317_),
    .Y(_11611_));
 sky130_fd_sc_hd__a31oi_4 _17128_ (.A1(net3599),
    .A2(_10964_),
    .A3(_11610_),
    .B1(_11611_),
    .Y(_11612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_788 ();
 sky130_fd_sc_hd__nor2_1 _17130_ (.A(net3491),
    .B(_11612_),
    .Y(_11614_));
 sky130_fd_sc_hd__a21oi_1 _17131_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(_11580_),
    .B1(_11614_),
    .Y(_11615_));
 sky130_fd_sc_hd__o21ai_0 _17132_ (.A1(_11147_),
    .A2(_11598_),
    .B1(_11615_),
    .Y(_00045_));
 sky130_fd_sc_hd__and3_1 _17133_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .C(_11590_),
    .X(_11616_));
 sky130_fd_sc_hd__nand2_1 _17134_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .B(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__nor3_1 _17135_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .B(_11574_),
    .C(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__a21oi_1 _17136_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(_11617_),
    .B1(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__a222oi_1 _17137_ (.A1(\cs_registers_i.csr_mepc_o[4] ),
    .A2(net3538),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[4] ),
    .C1(\cs_registers_i.csr_depc_o[4] ),
    .C2(_11221_),
    .Y(_11620_));
 sky130_fd_sc_hd__a22oi_1 _17138_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1860] ),
    .Y(_11621_));
 sky130_fd_sc_hd__a22oi_1 _17139_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1892] ),
    .Y(_11622_));
 sky130_fd_sc_hd__o22ai_1 _17140_ (.A1(_11130_),
    .A2(_11621_),
    .B1(_11622_),
    .B2(_11089_),
    .Y(_11623_));
 sky130_fd_sc_hd__nand2_2 _17141_ (.A(_11085_),
    .B(_11623_),
    .Y(_11624_));
 sky130_fd_sc_hd__a21oi_1 _17142_ (.A1(\cs_registers_i.mcause_q[4] ),
    .A2(_10613_),
    .B1(net3551),
    .Y(_11625_));
 sky130_fd_sc_hd__a22oi_1 _17143_ (.A1(\cs_registers_i.mscratch_q[4] ),
    .A2(net3540),
    .B1(net3552),
    .B2(net88),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(_11625_),
    .B(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__a221oi_1 _17145_ (.A1(\cs_registers_i.dscratch1_q[4] ),
    .A2(_11227_),
    .B1(_11228_),
    .B2(\cs_registers_i.dscratch0_q[4] ),
    .C1(_11627_),
    .Y(_11628_));
 sky130_fd_sc_hd__and3_4 _17146_ (.A(_11620_),
    .B(_11624_),
    .C(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__nand2_2 _17147_ (.A(net3594),
    .B(_10964_),
    .Y(_11630_));
 sky130_fd_sc_hd__o22ai_4 _17148_ (.A1(net3594),
    .A2(_11317_),
    .B1(_11629_),
    .B2(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__a22oi_1 _17149_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(_11580_),
    .B1(_11631_),
    .B2(_11579_),
    .Y(_11632_));
 sky130_fd_sc_hd__o21ai_0 _17150_ (.A1(_11147_),
    .A2(_11619_),
    .B1(_11632_),
    .Y(_00046_));
 sky130_fd_sc_hd__and2_0 _17151_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .B(_11616_),
    .X(_11633_));
 sky130_fd_sc_hd__nand2_1 _17152_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .B(_11633_),
    .Y(_11634_));
 sky130_fd_sc_hd__nor3_1 _17153_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .B(_11574_),
    .C(_11634_),
    .Y(_11635_));
 sky130_fd_sc_hd__a21oi_1 _17154_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_11634_),
    .B1(_11635_),
    .Y(_11636_));
 sky130_fd_sc_hd__a221o_4 _17155_ (.A1(\cs_registers_i.csr_mepc_o[5] ),
    .A2(net3538),
    .B1(_11057_),
    .B2(\cs_registers_i.dscratch0_q[5] ),
    .C1(_11052_),
    .X(_11637_));
 sky130_fd_sc_hd__a22oi_2 _17156_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1893] ),
    .Y(_11638_));
 sky130_fd_sc_hd__a22oi_1 _17157_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1861] ),
    .Y(_11639_));
 sky130_fd_sc_hd__o22ai_2 _17158_ (.A1(_11089_),
    .A2(_11638_),
    .B1(_11639_),
    .B2(_11130_),
    .Y(_11640_));
 sky130_fd_sc_hd__nand2_2 _17159_ (.A(_10993_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__a22oi_1 _17160_ (.A1(net89),
    .A2(_11070_),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[5] ),
    .Y(_11642_));
 sky130_fd_sc_hd__a22oi_2 _17161_ (.A1(\cs_registers_i.mtval_q[5] ),
    .A2(net3539),
    .B1(net3566),
    .B2(\cs_registers_i.csr_depc_o[5] ),
    .Y(_11643_));
 sky130_fd_sc_hd__nand3_2 _17162_ (.A(_11641_),
    .B(_11642_),
    .C(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__a211oi_4 _17163_ (.A1(\cs_registers_i.dscratch1_q[5] ),
    .A2(_11059_),
    .B1(_11637_),
    .C1(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__nor3_1 _17164_ (.A(net3600),
    .B(_10991_),
    .C(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__a21oi_4 _17165_ (.A1(net3600),
    .A2(_10965_),
    .B1(_11646_),
    .Y(_11647_));
 sky130_fd_sc_hd__nor2_1 _17166_ (.A(net3491),
    .B(_11647_),
    .Y(_11648_));
 sky130_fd_sc_hd__a21oi_1 _17167_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_11580_),
    .B1(_11648_),
    .Y(_11649_));
 sky130_fd_sc_hd__o21ai_0 _17168_ (.A1(_11147_),
    .A2(_11636_),
    .B1(_11649_),
    .Y(_00047_));
 sky130_fd_sc_hd__nand3_1 _17169_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .C(_11633_),
    .Y(_11650_));
 sky130_fd_sc_hd__nor3_1 _17170_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .B(_11574_),
    .C(_11650_),
    .Y(_11651_));
 sky130_fd_sc_hd__a21oi_1 _17171_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(_11650_),
    .B1(_11651_),
    .Y(_11652_));
 sky130_fd_sc_hd__a21oi_2 _17172_ (.A1(\cs_registers_i.dcsr_q[6] ),
    .A2(_11063_),
    .B1(_11052_),
    .Y(_11653_));
 sky130_fd_sc_hd__a22oi_1 _17173_ (.A1(net90),
    .A2(net3546),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[6] ),
    .Y(_11654_));
 sky130_fd_sc_hd__nand2_4 _17174_ (.A(_11653_),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__a221oi_2 _17175_ (.A1(\cs_registers_i.dscratch0_q[6] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[6] ),
    .C1(_11655_),
    .Y(_11656_));
 sky130_fd_sc_hd__a22oi_1 _17176_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1862] ),
    .Y(_11657_));
 sky130_fd_sc_hd__a22oi_2 _17177_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1894] ),
    .Y(_11658_));
 sky130_fd_sc_hd__o22ai_1 _17178_ (.A1(_11130_),
    .A2(_11657_),
    .B1(_11658_),
    .B2(_11089_),
    .Y(_11659_));
 sky130_fd_sc_hd__nand2_2 _17179_ (.A(_10993_),
    .B(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__a222oi_1 _17180_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(net3538),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[6] ),
    .C1(\cs_registers_i.csr_depc_o[6] ),
    .C2(net3566),
    .Y(_11661_));
 sky130_fd_sc_hd__and3_4 _17181_ (.A(_11656_),
    .B(_11660_),
    .C(net3526),
    .X(_11662_));
 sky130_fd_sc_hd__nor3_1 _17182_ (.A(net3601),
    .B(_10991_),
    .C(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__a21oi_4 _17183_ (.A1(net3601),
    .A2(_10965_),
    .B1(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(net3491),
    .B(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__a21oi_1 _17185_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(_11580_),
    .B1(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__o21ai_0 _17186_ (.A1(_11147_),
    .A2(_11652_),
    .B1(_11666_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _17187_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .Y(_11667_));
 sky130_fd_sc_hd__nand4_1 _17188_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .D(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .Y(_11668_));
 sky130_fd_sc_hd__nor2_2 _17189_ (.A(_11667_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__nand2_1 _17190_ (.A(_11590_),
    .B(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__nor3_1 _17191_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .B(_11574_),
    .C(_11670_),
    .Y(_11671_));
 sky130_fd_sc_hd__a21oi_1 _17192_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(_11670_),
    .B1(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__a221o_4 _17193_ (.A1(\cs_registers_i.mscratch_q[7] ),
    .A2(net3540),
    .B1(net3548),
    .B2(\cs_registers_i.dscratch0_q[7] ),
    .C1(_11052_),
    .X(_11673_));
 sky130_fd_sc_hd__a22oi_1 _17194_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1895] ),
    .Y(_11674_));
 sky130_fd_sc_hd__a22oi_1 _17195_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1863] ),
    .Y(_11675_));
 sky130_fd_sc_hd__o22ai_2 _17196_ (.A1(_11089_),
    .A2(_11674_),
    .B1(_11675_),
    .B2(_11130_),
    .Y(_11676_));
 sky130_fd_sc_hd__nand2_4 _17197_ (.A(_10993_),
    .B(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__a22o_4 _17198_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_11063_),
    .B1(_11076_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .X(_11678_));
 sky130_fd_sc_hd__a221oi_1 _17199_ (.A1(net147),
    .A2(_11104_),
    .B1(_10625_),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .C1(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__a22oi_1 _17200_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(_11098_),
    .B1(_10595_),
    .B2(\cs_registers_i.mstatus_q[4] ),
    .Y(_11680_));
 sky130_fd_sc_hd__a22oi_1 _17201_ (.A1(net91),
    .A2(net3546),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[7] ),
    .Y(_11681_));
 sky130_fd_sc_hd__nand4_1 _17202_ (.A(_11677_),
    .B(_11679_),
    .C(_11680_),
    .D(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__a211oi_4 _17203_ (.A1(\cs_registers_i.dscratch1_q[7] ),
    .A2(_11059_),
    .B1(_11673_),
    .C1(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__nor3_1 _17204_ (.A(_08810_),
    .B(_10991_),
    .C(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__a21oi_4 _17205_ (.A1(_08810_),
    .A2(_10965_),
    .B1(_11684_),
    .Y(_11685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_787 ();
 sky130_fd_sc_hd__nor2_1 _17207_ (.A(net3491),
    .B(net3478),
    .Y(_11687_));
 sky130_fd_sc_hd__a21oi_1 _17208_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(_11580_),
    .B1(_11687_),
    .Y(_11688_));
 sky130_fd_sc_hd__o21ai_0 _17209_ (.A1(_11147_),
    .A2(_11672_),
    .B1(_11688_),
    .Y(_00049_));
 sky130_fd_sc_hd__nand3_1 _17210_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .Y(_11689_));
 sky130_fd_sc_hd__o21ai_0 _17211_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_11689_),
    .B1(_11087_),
    .Y(_11690_));
 sky130_fd_sc_hd__a21oi_1 _17212_ (.A1(_11240_),
    .A2(_11690_),
    .B1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .Y(_11691_));
 sky130_fd_sc_hd__and3_1 _17213_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .B(_11113_),
    .C(_11150_),
    .X(_11692_));
 sky130_fd_sc_hd__a211oi_1 _17214_ (.A1(_11120_),
    .A2(_11612_),
    .B1(_11691_),
    .C1(_11692_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand3_1 _17215_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .B(_11590_),
    .C(_11669_),
    .Y(_11693_));
 sky130_fd_sc_hd__nor3_1 _17216_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .B(_11574_),
    .C(_11693_),
    .Y(_11694_));
 sky130_fd_sc_hd__a21oi_1 _17217_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(_11693_),
    .B1(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__a22oi_2 _17218_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1896] ),
    .Y(_11696_));
 sky130_fd_sc_hd__a22oi_1 _17219_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1864] ),
    .Y(_11697_));
 sky130_fd_sc_hd__o22ai_4 _17220_ (.A1(_11089_),
    .A2(_11696_),
    .B1(_11697_),
    .B2(_11130_),
    .Y(_11698_));
 sky130_fd_sc_hd__a22o_1 _17221_ (.A1(\cs_registers_i.csr_mtvec_o[8] ),
    .A2(net3550),
    .B1(_11342_),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .X(_11699_));
 sky130_fd_sc_hd__a221o_4 _17222_ (.A1(\cs_registers_i.mscratch_q[8] ),
    .A2(net3540),
    .B1(net3539),
    .B2(\cs_registers_i.mtval_q[8] ),
    .C1(_11699_),
    .X(_11700_));
 sky130_fd_sc_hd__nand2_1 _17223_ (.A(net92),
    .B(net3552),
    .Y(_11701_));
 sky130_fd_sc_hd__a22oi_2 _17224_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(net3538),
    .B1(_11221_),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .Y(_11702_));
 sky130_fd_sc_hd__a22oi_1 _17225_ (.A1(\cs_registers_i.dscratch1_q[8] ),
    .A2(_11227_),
    .B1(_11228_),
    .B2(\cs_registers_i.dscratch0_q[8] ),
    .Y(_11703_));
 sky130_fd_sc_hd__nand4_1 _17226_ (.A(_10608_),
    .B(_11701_),
    .C(_11702_),
    .D(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__a211oi_4 _17227_ (.A1(_11085_),
    .A2(_11698_),
    .B1(_11700_),
    .C1(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__nor3_1 _17228_ (.A(net3615),
    .B(_10991_),
    .C(_11705_),
    .Y(_11706_));
 sky130_fd_sc_hd__a21oi_4 _17229_ (.A1(net3615),
    .A2(_10965_),
    .B1(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_786 ();
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(net3491),
    .B(_11707_),
    .Y(_11709_));
 sky130_fd_sc_hd__a21oi_1 _17232_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(_11580_),
    .B1(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__o21ai_0 _17233_ (.A1(_11147_),
    .A2(_11695_),
    .B1(_11710_),
    .Y(_00051_));
 sky130_fd_sc_hd__nand3_1 _17234_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .C(_11669_),
    .Y(_11711_));
 sky130_fd_sc_hd__or2_0 _17235_ (.A(_11585_),
    .B(_11711_),
    .X(_11712_));
 sky130_fd_sc_hd__nor3_1 _17236_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .B(_11574_),
    .C(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__a21oi_1 _17237_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(_11712_),
    .B1(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__a21oi_1 _17238_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(net3539),
    .B1(_11052_),
    .Y(_11715_));
 sky130_fd_sc_hd__a22oi_2 _17239_ (.A1(net93),
    .A2(net3546),
    .B1(net3538),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .Y(_11716_));
 sky130_fd_sc_hd__nand2_4 _17240_ (.A(_11715_),
    .B(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__a221oi_1 _17241_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(_11057_),
    .B1(_11059_),
    .B2(\cs_registers_i.dscratch1_q[9] ),
    .C1(_11717_),
    .Y(_11718_));
 sky130_fd_sc_hd__a22oi_1 _17242_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1865] ),
    .Y(_11719_));
 sky130_fd_sc_hd__a22oi_2 _17243_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(net3581),
    .B1(_10610_),
    .B2(\cs_registers_i.mhpmcounter[1897] ),
    .Y(_11720_));
 sky130_fd_sc_hd__o22ai_2 _17244_ (.A1(_11130_),
    .A2(_11719_),
    .B1(_11720_),
    .B2(_11089_),
    .Y(_11721_));
 sky130_fd_sc_hd__nand2_2 _17245_ (.A(_10993_),
    .B(_11721_),
    .Y(_11722_));
 sky130_fd_sc_hd__a222oi_1 _17246_ (.A1(\cs_registers_i.csr_mtvec_o[9] ),
    .A2(net3550),
    .B1(net3540),
    .B2(\cs_registers_i.mscratch_q[9] ),
    .C1(net3566),
    .C2(\cs_registers_i.csr_depc_o[9] ),
    .Y(_11723_));
 sky130_fd_sc_hd__and3_4 _17247_ (.A(_11718_),
    .B(_11722_),
    .C(net3525),
    .X(_11724_));
 sky130_fd_sc_hd__nor3_1 _17248_ (.A(net3617),
    .B(_10991_),
    .C(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__a21oi_4 _17249_ (.A1(net3617),
    .A2(_10965_),
    .B1(_11725_),
    .Y(_11726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_785 ();
 sky130_fd_sc_hd__nor2_1 _17251_ (.A(net3491),
    .B(_11726_),
    .Y(_11728_));
 sky130_fd_sc_hd__a21oi_1 _17252_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(_11580_),
    .B1(_11728_),
    .Y(_11729_));
 sky130_fd_sc_hd__o21ai_0 _17253_ (.A1(_11147_),
    .A2(_11714_),
    .B1(_11729_),
    .Y(_00052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_784 ();
 sky130_fd_sc_hd__nor2_1 _17255_ (.A(_11585_),
    .B(_11711_),
    .Y(_11731_));
 sky130_fd_sc_hd__nand2_1 _17256_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .B(_11731_),
    .Y(_11732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_783 ();
 sky130_fd_sc_hd__nor3_1 _17258_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .B(_11574_),
    .C(_11732_),
    .Y(_11734_));
 sky130_fd_sc_hd__a21oi_1 _17259_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(_11732_),
    .B1(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__nor2_1 _17260_ (.A(_11145_),
    .B(net3491),
    .Y(_11736_));
 sky130_fd_sc_hd__a21oi_1 _17261_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(_11580_),
    .B1(_11736_),
    .Y(_11737_));
 sky130_fd_sc_hd__o21ai_0 _17262_ (.A1(_11147_),
    .A2(_11735_),
    .B1(_11737_),
    .Y(_00053_));
 sky130_fd_sc_hd__nand3_1 _17263_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .Y(_11738_));
 sky130_fd_sc_hd__or3_4 _17264_ (.A(_11572_),
    .B(_11711_),
    .C(_11738_),
    .X(_11739_));
 sky130_fd_sc_hd__nor3_1 _17265_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .B(_11574_),
    .C(_11739_),
    .Y(_11740_));
 sky130_fd_sc_hd__a21oi_1 _17266_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_11739_),
    .B1(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_782 ();
 sky130_fd_sc_hd__nor2_1 _17268_ (.A(_11177_),
    .B(net3491),
    .Y(_11743_));
 sky130_fd_sc_hd__a21oi_1 _17269_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_11580_),
    .B1(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__o21ai_0 _17270_ (.A1(net3484),
    .A2(_11741_),
    .B1(_11744_),
    .Y(_00054_));
 sky130_fd_sc_hd__clkinv_1 _17271_ (.A(_11739_),
    .Y(_11745_));
 sky130_fd_sc_hd__nand2_2 _17272_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .B(_11745_),
    .Y(_11746_));
 sky130_fd_sc_hd__nor3_1 _17273_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .B(_11574_),
    .C(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__a21oi_1 _17274_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_11746_),
    .B1(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__nor2_1 _17275_ (.A(_11197_),
    .B(net3491),
    .Y(_11749_));
 sky130_fd_sc_hd__a21oi_1 _17276_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_11580_),
    .B1(_11749_),
    .Y(_11750_));
 sky130_fd_sc_hd__o21ai_0 _17277_ (.A1(net3484),
    .A2(_11748_),
    .B1(_11750_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand3_1 _17278_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .C(_11745_),
    .Y(_11751_));
 sky130_fd_sc_hd__nor3_1 _17279_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .B(_11574_),
    .C(_11751_),
    .Y(_11752_));
 sky130_fd_sc_hd__a21oi_1 _17280_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(_11751_),
    .B1(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__nor2_1 _17281_ (.A(_11214_),
    .B(net3491),
    .Y(_11754_));
 sky130_fd_sc_hd__a21oi_1 _17282_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(_11580_),
    .B1(_11754_),
    .Y(_11755_));
 sky130_fd_sc_hd__o21ai_0 _17283_ (.A1(net3484),
    .A2(_11753_),
    .B1(_11755_),
    .Y(_00056_));
 sky130_fd_sc_hd__and3_4 _17284_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .C(_11745_),
    .X(_11756_));
 sky130_fd_sc_hd__nand2_1 _17285_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .B(_11756_),
    .Y(_11757_));
 sky130_fd_sc_hd__nor3_1 _17286_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .B(_11574_),
    .C(_11757_),
    .Y(_11758_));
 sky130_fd_sc_hd__a21oi_1 _17287_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_11757_),
    .B1(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__nor2_1 _17288_ (.A(_11235_),
    .B(net3491),
    .Y(_11760_));
 sky130_fd_sc_hd__a21oi_1 _17289_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_11580_),
    .B1(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__o21ai_0 _17290_ (.A1(net3484),
    .A2(_11759_),
    .B1(_11761_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand3_1 _17291_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .C(_11756_),
    .Y(_11762_));
 sky130_fd_sc_hd__nor3_1 _17292_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .B(_11574_),
    .C(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__a21oi_1 _17293_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(_11762_),
    .B1(_11763_),
    .Y(_11764_));
 sky130_fd_sc_hd__nor2_1 _17294_ (.A(_11255_),
    .B(net3491),
    .Y(_11765_));
 sky130_fd_sc_hd__a21oi_1 _17295_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(_11580_),
    .B1(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__o21ai_0 _17296_ (.A1(net3484),
    .A2(_11764_),
    .B1(_11766_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand4_1 _17297_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .D(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .Y(_11767_));
 sky130_fd_sc_hd__nor2_2 _17298_ (.A(_11746_),
    .B(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__inv_1 _17299_ (.A(_11768_),
    .Y(_11769_));
 sky130_fd_sc_hd__nor3_1 _17300_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .B(_11574_),
    .C(_11769_),
    .Y(_11770_));
 sky130_fd_sc_hd__a21oi_1 _17301_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(_11769_),
    .B1(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__nor2_1 _17302_ (.A(_11270_),
    .B(net3491),
    .Y(_11772_));
 sky130_fd_sc_hd__a21oi_1 _17303_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(_11580_),
    .B1(_11772_),
    .Y(_11773_));
 sky130_fd_sc_hd__o21ai_0 _17304_ (.A1(net3484),
    .A2(_11771_),
    .B1(_11773_),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _17305_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .B(_11768_),
    .Y(_11774_));
 sky130_fd_sc_hd__nor3_1 _17306_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .B(_11574_),
    .C(_11774_),
    .Y(_11775_));
 sky130_fd_sc_hd__a21oi_1 _17307_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(_11774_),
    .B1(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_781 ();
 sky130_fd_sc_hd__nor2_1 _17309_ (.A(_11294_),
    .B(net3491),
    .Y(_11778_));
 sky130_fd_sc_hd__a21oi_1 _17310_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(_11580_),
    .B1(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__o21ai_0 _17311_ (.A1(net3484),
    .A2(_11776_),
    .B1(_11779_),
    .Y(_00060_));
 sky130_fd_sc_hd__o22a_4 _17312_ (.A1(net3594),
    .A2(_11317_),
    .B1(_11629_),
    .B2(_11630_),
    .X(_11780_));
 sky130_fd_sc_hd__nor3_1 _17313_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .B(_11115_),
    .C(_11692_),
    .Y(_11781_));
 sky130_fd_sc_hd__nor3_2 _17314_ (.A(\cs_registers_i.mcountinhibit_q[0] ),
    .B(net3484),
    .C(_11151_),
    .Y(_11782_));
 sky130_fd_sc_hd__a211oi_1 _17315_ (.A1(_11115_),
    .A2(_11780_),
    .B1(_11781_),
    .C1(_11782_),
    .Y(_00061_));
 sky130_fd_sc_hd__and2_4 _17316_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .B(_11768_),
    .X(_11783_));
 sky130_fd_sc_hd__nand2_1 _17317_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .B(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__nor3_1 _17318_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .B(_11574_),
    .C(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__a21oi_1 _17319_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(_11784_),
    .B1(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__nor2_1 _17320_ (.A(_11319_),
    .B(net3491),
    .Y(_11787_));
 sky130_fd_sc_hd__a21oi_1 _17321_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(_11580_),
    .B1(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__o21ai_0 _17322_ (.A1(net3484),
    .A2(_11786_),
    .B1(_11788_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand3_1 _17323_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .C(_11783_),
    .Y(_11789_));
 sky130_fd_sc_hd__nor3_1 _17324_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .B(_11574_),
    .C(_11789_),
    .Y(_11790_));
 sky130_fd_sc_hd__a21oi_1 _17325_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(_11789_),
    .B1(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__nor2_1 _17326_ (.A(_11333_),
    .B(net3491),
    .Y(_11792_));
 sky130_fd_sc_hd__a21oi_1 _17327_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(_11580_),
    .B1(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__o21ai_0 _17328_ (.A1(net3484),
    .A2(_11791_),
    .B1(_11793_),
    .Y(_00063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_780 ();
 sky130_fd_sc_hd__and3_4 _17330_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .C(_11783_),
    .X(_11795_));
 sky130_fd_sc_hd__nand2_1 _17331_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .B(_11795_),
    .Y(_11796_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_779 ();
 sky130_fd_sc_hd__nor3_1 _17333_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .B(_11574_),
    .C(_11796_),
    .Y(_11798_));
 sky130_fd_sc_hd__a21oi_1 _17334_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(_11796_),
    .B1(_11798_),
    .Y(_11799_));
 sky130_fd_sc_hd__nor2_1 _17335_ (.A(_11369_),
    .B(net3491),
    .Y(_11800_));
 sky130_fd_sc_hd__a21oi_1 _17336_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(_11580_),
    .B1(_11800_),
    .Y(_11801_));
 sky130_fd_sc_hd__o21ai_0 _17337_ (.A1(net3484),
    .A2(_11799_),
    .B1(_11801_),
    .Y(_00064_));
 sky130_fd_sc_hd__and2_4 _17338_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .B(_11795_),
    .X(_11802_));
 sky130_fd_sc_hd__nand2_1 _17339_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .B(_11802_),
    .Y(_11803_));
 sky130_fd_sc_hd__nor3_1 _17340_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .B(_11574_),
    .C(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__a21oi_1 _17341_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(_11803_),
    .B1(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_778 ();
 sky130_fd_sc_hd__nor2_1 _17343_ (.A(net3494),
    .B(net3491),
    .Y(_11807_));
 sky130_fd_sc_hd__a21oi_1 _17344_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(_11580_),
    .B1(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__o21ai_0 _17345_ (.A1(net3484),
    .A2(_11805_),
    .B1(_11808_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand3_1 _17346_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .C(_11802_),
    .Y(_11809_));
 sky130_fd_sc_hd__nor3_1 _17347_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .B(_11574_),
    .C(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__a21oi_1 _17348_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_11809_),
    .B1(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(net3493),
    .B(net3491),
    .Y(_11812_));
 sky130_fd_sc_hd__a21oi_1 _17350_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_11580_),
    .B1(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__o21ai_0 _17351_ (.A1(net3484),
    .A2(_11811_),
    .B1(_11813_),
    .Y(_00066_));
 sky130_fd_sc_hd__and3_1 _17352_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .C(_11802_),
    .X(_11814_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .B(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__nor3_1 _17354_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .B(_11574_),
    .C(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__a21oi_1 _17355_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(_11815_),
    .B1(_11816_),
    .Y(_11817_));
 sky130_fd_sc_hd__nor2_1 _17356_ (.A(net3492),
    .B(net3491),
    .Y(_11818_));
 sky130_fd_sc_hd__a21oi_1 _17357_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(_11580_),
    .B1(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__o21ai_0 _17358_ (.A1(net3484),
    .A2(_11817_),
    .B1(_11819_),
    .Y(_00067_));
 sky130_fd_sc_hd__and2_4 _17359_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .B(_11814_),
    .X(_11820_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .B(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__nor3_1 _17361_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .B(_11574_),
    .C(_11821_),
    .Y(_11822_));
 sky130_fd_sc_hd__a21oi_1 _17362_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(_11821_),
    .B1(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__nor2_1 _17363_ (.A(net3483),
    .B(net3491),
    .Y(_11824_));
 sky130_fd_sc_hd__a21oi_1 _17364_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(_11580_),
    .B1(_11824_),
    .Y(_11825_));
 sky130_fd_sc_hd__o21ai_0 _17365_ (.A1(net3484),
    .A2(_11823_),
    .B1(_11825_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand3_1 _17366_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .C(_11820_),
    .Y(_11826_));
 sky130_fd_sc_hd__nor3_1 _17367_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .B(_11574_),
    .C(_11826_),
    .Y(_11827_));
 sky130_fd_sc_hd__a21oi_1 _17368_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(_11826_),
    .B1(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__nor2_1 _17369_ (.A(_11457_),
    .B(net3491),
    .Y(_11829_));
 sky130_fd_sc_hd__a21oi_1 _17370_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(_11580_),
    .B1(_11829_),
    .Y(_11830_));
 sky130_fd_sc_hd__o21ai_0 _17371_ (.A1(net3484),
    .A2(_11828_),
    .B1(_11830_),
    .Y(_00069_));
 sky130_fd_sc_hd__and3_4 _17372_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .C(_11820_),
    .X(_11831_));
 sky130_fd_sc_hd__nand2_1 _17373_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .B(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__nor3_1 _17374_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .B(_11574_),
    .C(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__a21oi_1 _17375_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(_11832_),
    .B1(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__nor2_1 _17376_ (.A(net3482),
    .B(net3491),
    .Y(_11835_));
 sky130_fd_sc_hd__a21oi_1 _17377_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(_11580_),
    .B1(_11835_),
    .Y(_11836_));
 sky130_fd_sc_hd__o21ai_0 _17378_ (.A1(net3484),
    .A2(_11834_),
    .B1(_11836_),
    .Y(_00070_));
 sky130_fd_sc_hd__and2_4 _17379_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .B(_11831_),
    .X(_11837_));
 sky130_fd_sc_hd__nand2_1 _17380_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .B(_11837_),
    .Y(_11838_));
 sky130_fd_sc_hd__nor3_1 _17381_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .B(_11574_),
    .C(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__a21oi_1 _17382_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(_11838_),
    .B1(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__nor2_1 _17383_ (.A(net3481),
    .B(net3491),
    .Y(_11841_));
 sky130_fd_sc_hd__a21oi_1 _17384_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(_11580_),
    .B1(_11841_),
    .Y(_11842_));
 sky130_fd_sc_hd__o21ai_0 _17385_ (.A1(net3484),
    .A2(_11840_),
    .B1(_11842_),
    .Y(_00071_));
 sky130_fd_sc_hd__a22oi_1 _17386_ (.A1(_11115_),
    .A2(_11647_),
    .B1(_11782_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .Y(_11843_));
 sky130_fd_sc_hd__o31a_1 _17387_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .A2(_11115_),
    .A3(_11782_),
    .B1(_11843_),
    .X(_00072_));
 sky130_fd_sc_hd__nand3_1 _17388_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .C(_11837_),
    .Y(_11844_));
 sky130_fd_sc_hd__nor3_1 _17389_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .B(_11574_),
    .C(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__a21oi_1 _17390_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(_11844_),
    .B1(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__nor2_1 _17391_ (.A(net3480),
    .B(net3491),
    .Y(_11847_));
 sky130_fd_sc_hd__a21oi_1 _17392_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(_11580_),
    .B1(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21ai_0 _17393_ (.A1(net3484),
    .A2(_11846_),
    .B1(_11848_),
    .Y(_00073_));
 sky130_fd_sc_hd__and3_4 _17394_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .C(_11837_),
    .X(_11849_));
 sky130_fd_sc_hd__nand2_1 _17395_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .B(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__nor3_1 _17396_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .B(_11574_),
    .C(_11850_),
    .Y(_11851_));
 sky130_fd_sc_hd__a21oi_1 _17397_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(_11850_),
    .B1(_11851_),
    .Y(_11852_));
 sky130_fd_sc_hd__nor2_1 _17398_ (.A(net3479),
    .B(net3491),
    .Y(_11853_));
 sky130_fd_sc_hd__a21oi_1 _17399_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(_11580_),
    .B1(_11853_),
    .Y(_11854_));
 sky130_fd_sc_hd__o21ai_0 _17400_ (.A1(net3484),
    .A2(_11852_),
    .B1(_11854_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand3_1 _17401_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .C(_11849_),
    .Y(_11855_));
 sky130_fd_sc_hd__nor3_1 _17402_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .B(_11574_),
    .C(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__a21oi_1 _17403_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(_11855_),
    .B1(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__nor2_1 _17404_ (.A(_11550_),
    .B(net3491),
    .Y(_11858_));
 sky130_fd_sc_hd__a21oi_1 _17405_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(_11580_),
    .B1(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__o21ai_0 _17406_ (.A1(net3484),
    .A2(_11857_),
    .B1(_11859_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand4_1 _17407_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .D(_11849_),
    .Y(_11860_));
 sky130_fd_sc_hd__nor3_1 _17408_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .B(_11574_),
    .C(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__a21oi_1 _17409_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(_11860_),
    .B1(_11861_),
    .Y(_11862_));
 sky130_fd_sc_hd__nor2_1 _17410_ (.A(_11565_),
    .B(net3491),
    .Y(_11863_));
 sky130_fd_sc_hd__a21oi_1 _17411_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(_11580_),
    .B1(_11863_),
    .Y(_11864_));
 sky130_fd_sc_hd__o21ai_0 _17412_ (.A1(net3484),
    .A2(_11862_),
    .B1(_11864_),
    .Y(_00076_));
 sky130_fd_sc_hd__a211oi_1 _17413_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .A2(_11782_),
    .B1(_11120_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .Y(_11865_));
 sky130_fd_sc_hd__and3_1 _17414_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .C(_11782_),
    .X(_11866_));
 sky130_fd_sc_hd__a211oi_1 _17415_ (.A1(_11115_),
    .A2(_11664_),
    .B1(_11865_),
    .C1(_11866_),
    .Y(_00077_));
 sky130_fd_sc_hd__o21ai_0 _17416_ (.A1(net3484),
    .A2(_11152_),
    .B1(_11240_),
    .Y(_11867_));
 sky130_fd_sc_hd__nand2_1 _17417_ (.A(_11087_),
    .B(_11152_),
    .Y(_11868_));
 sky130_fd_sc_hd__o22ai_1 _17418_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(_11868_),
    .B1(net3478),
    .B2(_11202_),
    .Y(_11869_));
 sky130_fd_sc_hd__a21o_1 _17419_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(_11867_),
    .B1(_11869_),
    .X(_00078_));
 sky130_fd_sc_hd__a311oi_1 _17420_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(_11087_),
    .A3(_11152_),
    .B1(_11115_),
    .C1(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .Y(_11870_));
 sky130_fd_sc_hd__a211oi_1 _17421_ (.A1(_11115_),
    .A2(_11707_),
    .B1(_11870_),
    .C1(_11154_),
    .Y(_00079_));
 sky130_fd_sc_hd__inv_1 _17422_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .Y(_11871_));
 sky130_fd_sc_hd__a21oi_1 _17423_ (.A1(_11087_),
    .A2(_11153_),
    .B1(_11091_),
    .Y(_11872_));
 sky130_fd_sc_hd__nor2_1 _17424_ (.A(_11202_),
    .B(_11726_),
    .Y(_11873_));
 sky130_fd_sc_hd__a21oi_1 _17425_ (.A1(_11871_),
    .A2(_11154_),
    .B1(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__o21ai_0 _17426_ (.A1(_11871_),
    .A2(_11872_),
    .B1(_11874_),
    .Y(_00080_));
 sky130_fd_sc_hd__nor2_4 _17427_ (.A(_11002_),
    .B(_11004_),
    .Y(_11875_));
 sky130_fd_sc_hd__inv_1 _17428_ (.A(_10999_),
    .Y(_11876_));
 sky130_fd_sc_hd__o21ai_0 _17429_ (.A1(_11876_),
    .A2(_10554_),
    .B1(_11019_),
    .Y(_11877_));
 sky130_fd_sc_hd__a21oi_1 _17430_ (.A1(_10553_),
    .A2(_11877_),
    .B1(_11364_),
    .Y(_11878_));
 sky130_fd_sc_hd__nor2_1 _17431_ (.A(_11036_),
    .B(_10585_),
    .Y(_11879_));
 sky130_fd_sc_hd__or4_4 _17432_ (.A(_11028_),
    .B(_11029_),
    .C(_11879_),
    .D(_11035_),
    .X(_11880_));
 sky130_fd_sc_hd__a2111oi_0 _17433_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11032_),
    .C1(_11312_),
    .D1(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__nor4_1 _17434_ (.A(_11017_),
    .B(_10587_),
    .C(_10616_),
    .D(_11094_),
    .Y(_11882_));
 sky130_fd_sc_hd__a2111oi_0 _17435_ (.A1(_10622_),
    .A2(_11882_),
    .B1(_11307_),
    .C1(_11033_),
    .D1(_11037_),
    .Y(_11883_));
 sky130_fd_sc_hd__nand4_1 _17436_ (.A(_11878_),
    .B(_11881_),
    .C(_11875_),
    .D(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__o2111a_4 _17437_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_11019_),
    .B1(_11884_),
    .C1(_10635_),
    .D1(_11110_),
    .X(_11885_));
 sky130_fd_sc_hd__nand2_2 _17438_ (.A(_10993_),
    .B(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__nor3_4 _17439_ (.A(_11875_),
    .B(_11009_),
    .C(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__nand2_8 _17440_ (.A(_11303_),
    .B(net3490),
    .Y(_11888_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_777 ();
 sky130_fd_sc_hd__nand2_8 _17442_ (.A(_10542_),
    .B(_10639_),
    .Y(_11890_));
 sky130_fd_sc_hd__nand3_1 _17443_ (.A(net3750),
    .B(net3785),
    .C(_10517_),
    .Y(_11891_));
 sky130_fd_sc_hd__nor2_1 _17444_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(\cs_registers_i.mcountinhibit_q[2] ),
    .Y(_11892_));
 sky130_fd_sc_hd__nand3_4 _17445_ (.A(_10655_),
    .B(_11891_),
    .C(_11892_),
    .Y(_11893_));
 sky130_fd_sc_hd__nor4_2 _17446_ (.A(net3449),
    .B(_11887_),
    .C(_11890_),
    .D(_11893_),
    .Y(_11894_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_775 ();
 sky130_fd_sc_hd__or4_4 _17449_ (.A(net3449),
    .B(_11887_),
    .C(_11890_),
    .D(_11893_),
    .X(_11897_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_774 ();
 sky130_fd_sc_hd__nand2_8 _17451_ (.A(_11888_),
    .B(_11897_),
    .Y(_11899_));
 sky130_fd_sc_hd__nand2_1 _17452_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(_11899_),
    .Y(_11900_));
 sky130_fd_sc_hd__o21ai_0 _17453_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(net3439),
    .B1(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__o21ai_0 _17454_ (.A1(_11042_),
    .A2(_11888_),
    .B1(_11901_),
    .Y(_00081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_773 ();
 sky130_fd_sc_hd__and4_4 _17456_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .C(\cs_registers_i.mhpmcounter[1858] ),
    .D(\cs_registers_i.mhpmcounter[1859] ),
    .X(_11903_));
 sky130_fd_sc_hd__and3_4 _17457_ (.A(\cs_registers_i.mhpmcounter[1860] ),
    .B(\cs_registers_i.mhpmcounter[1861] ),
    .C(_11903_),
    .X(_11904_));
 sky130_fd_sc_hd__and3_4 _17458_ (.A(\cs_registers_i.mhpmcounter[1862] ),
    .B(\cs_registers_i.mhpmcounter[1863] ),
    .C(_11904_),
    .X(_11905_));
 sky130_fd_sc_hd__nand4_1 _17459_ (.A(\cs_registers_i.mhpmcounter[1864] ),
    .B(\cs_registers_i.mhpmcounter[1865] ),
    .C(net3435),
    .D(_11905_),
    .Y(_11906_));
 sky130_fd_sc_hd__xnor2_1 _17460_ (.A(\cs_registers_i.mhpmcounter[1866] ),
    .B(_11906_),
    .Y(_11907_));
 sky130_fd_sc_hd__nand2_1 _17461_ (.A(_11888_),
    .B(_11907_),
    .Y(_11908_));
 sky130_fd_sc_hd__o21ai_0 _17462_ (.A1(_11145_),
    .A2(_11888_),
    .B1(_11908_),
    .Y(_00082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_771 ();
 sky130_fd_sc_hd__and2_4 _17465_ (.A(\cs_registers_i.mhpmcounter[1862] ),
    .B(_11904_),
    .X(_11911_));
 sky130_fd_sc_hd__nand2_2 _17466_ (.A(\cs_registers_i.mhpmcounter[1863] ),
    .B(_11911_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand3_2 _17467_ (.A(\cs_registers_i.mhpmcounter[1864] ),
    .B(\cs_registers_i.mhpmcounter[1865] ),
    .C(\cs_registers_i.mhpmcounter[1866] ),
    .Y(_11913_));
 sky130_fd_sc_hd__nor2_1 _17468_ (.A(_11912_),
    .B(_11913_),
    .Y(_11914_));
 sky130_fd_sc_hd__nand3b_1 _17469_ (.A_N(\cs_registers_i.mhpmcounter[1867] ),
    .B(net3435),
    .C(_11914_),
    .Y(_11915_));
 sky130_fd_sc_hd__or3_4 _17470_ (.A(_11875_),
    .B(_11009_),
    .C(_11886_),
    .X(_11916_));
 sky130_fd_sc_hd__nor2_2 _17471_ (.A(_11004_),
    .B(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__nor2_4 _17472_ (.A(_11917_),
    .B(net3435),
    .Y(_11918_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_769 ();
 sky130_fd_sc_hd__nor2_1 _17475_ (.A(net3434),
    .B(_11914_),
    .Y(_11921_));
 sky130_fd_sc_hd__o21ai_0 _17476_ (.A1(_11918_),
    .A2(_11921_),
    .B1(\cs_registers_i.mhpmcounter[1867] ),
    .Y(_11922_));
 sky130_fd_sc_hd__o211ai_1 _17477_ (.A1(_11177_),
    .A2(_11888_),
    .B1(_11915_),
    .C1(_11922_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _17478_ (.A(\cs_registers_i.mhpmcounter[1867] ),
    .B(_11914_),
    .Y(_11923_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_11897_),
    .B(_11923_),
    .Y(_11924_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_768 ();
 sky130_fd_sc_hd__nand2_1 _17481_ (.A(net3436),
    .B(_11923_),
    .Y(_11926_));
 sky130_fd_sc_hd__nand3_1 _17482_ (.A(\cs_registers_i.mhpmcounter[1868] ),
    .B(_11899_),
    .C(_11926_),
    .Y(_11927_));
 sky130_fd_sc_hd__o21ai_0 _17483_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(net3427),
    .B1(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__o21ai_0 _17484_ (.A1(_11197_),
    .A2(_11888_),
    .B1(_11928_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _17485_ (.A(\cs_registers_i.mhpmcounter[1868] ),
    .B(net3427),
    .Y(_11929_));
 sky130_fd_sc_hd__nor2_4 _17486_ (.A(_11303_),
    .B(net3435),
    .Y(_11930_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_766 ();
 sky130_fd_sc_hd__a21oi_1 _17489_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(_11924_),
    .B1(net3490),
    .Y(_11933_));
 sky130_fd_sc_hd__o21ai_0 _17490_ (.A1(_11930_),
    .A2(_11933_),
    .B1(\cs_registers_i.mhpmcounter[1869] ),
    .Y(_11934_));
 sky130_fd_sc_hd__o221ai_1 _17491_ (.A1(_11214_),
    .A2(_11888_),
    .B1(_11929_),
    .B2(\cs_registers_i.mhpmcounter[1869] ),
    .C1(_11934_),
    .Y(_00085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_765 ();
 sky130_fd_sc_hd__nand3_1 _17493_ (.A(\cs_registers_i.mhpmcounter[1868] ),
    .B(\cs_registers_i.mhpmcounter[1867] ),
    .C(\cs_registers_i.mhpmcounter[1869] ),
    .Y(_11936_));
 sky130_fd_sc_hd__nor3_2 _17494_ (.A(_11912_),
    .B(_11913_),
    .C(_11936_),
    .Y(_11937_));
 sky130_fd_sc_hd__o211a_1 _17495_ (.A1(net3434),
    .A2(_11937_),
    .B1(_11899_),
    .C1(\cs_registers_i.mhpmcounter[1870] ),
    .X(_11938_));
 sky130_fd_sc_hd__a21oi_1 _17496_ (.A1(net3437),
    .A2(_11937_),
    .B1(\cs_registers_i.mhpmcounter[1870] ),
    .Y(_11939_));
 sky130_fd_sc_hd__o22ai_1 _17497_ (.A1(_11235_),
    .A2(_11888_),
    .B1(_11938_),
    .B2(_11939_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand4b_1 _17498_ (.A_N(\cs_registers_i.mhpmcounter[1871] ),
    .B(net3437),
    .C(_11937_),
    .D(\cs_registers_i.mhpmcounter[1870] ),
    .Y(_11940_));
 sky130_fd_sc_hd__a21oi_1 _17499_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(_11937_),
    .B1(net3434),
    .Y(_11941_));
 sky130_fd_sc_hd__o21ai_0 _17500_ (.A1(_11918_),
    .A2(_11941_),
    .B1(\cs_registers_i.mhpmcounter[1871] ),
    .Y(_11942_));
 sky130_fd_sc_hd__o211ai_1 _17501_ (.A1(_11255_),
    .A2(_11888_),
    .B1(_11940_),
    .C1(_11942_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand4_1 _17502_ (.A(\cs_registers_i.mhpmcounter[1870] ),
    .B(\cs_registers_i.mhpmcounter[1871] ),
    .C(net3435),
    .D(_11937_),
    .Y(_11943_));
 sky130_fd_sc_hd__xnor2_1 _17503_ (.A(\cs_registers_i.mhpmcounter[1872] ),
    .B(_11943_),
    .Y(_11944_));
 sky130_fd_sc_hd__nand2_1 _17504_ (.A(_11888_),
    .B(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__o21ai_0 _17505_ (.A1(_11270_),
    .A2(_11888_),
    .B1(_11945_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand3_1 _17506_ (.A(\cs_registers_i.mhpmcounter[1870] ),
    .B(\cs_registers_i.mhpmcounter[1871] ),
    .C(\cs_registers_i.mhpmcounter[1872] ),
    .Y(_11946_));
 sky130_fd_sc_hd__nor3_1 _17507_ (.A(_11913_),
    .B(_11936_),
    .C(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__and3_1 _17508_ (.A(net3435),
    .B(_11905_),
    .C(_11947_),
    .X(_11948_));
 sky130_fd_sc_hd__o221ai_1 _17509_ (.A1(_11303_),
    .A2(net3435),
    .B1(_11948_),
    .B2(net3490),
    .C1(\cs_registers_i.mhpmcounter[1873] ),
    .Y(_11949_));
 sky130_fd_sc_hd__o21ai_0 _17510_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(_11948_),
    .B1(_11949_),
    .Y(_11950_));
 sky130_fd_sc_hd__o21ai_0 _17511_ (.A1(_11294_),
    .A2(_11888_),
    .B1(_11950_),
    .Y(_00089_));
 sky130_fd_sc_hd__and3_4 _17512_ (.A(\cs_registers_i.mhpmcounter[1873] ),
    .B(_11905_),
    .C(_11947_),
    .X(_11951_));
 sky130_fd_sc_hd__o211a_1 _17513_ (.A1(net3434),
    .A2(_11951_),
    .B1(_11899_),
    .C1(\cs_registers_i.mhpmcounter[1874] ),
    .X(_11952_));
 sky130_fd_sc_hd__a21oi_1 _17514_ (.A1(net3438),
    .A2(_11951_),
    .B1(\cs_registers_i.mhpmcounter[1874] ),
    .Y(_11953_));
 sky130_fd_sc_hd__o22ai_1 _17515_ (.A1(_11319_),
    .A2(_11888_),
    .B1(_11952_),
    .B2(_11953_),
    .Y(_00090_));
 sky130_fd_sc_hd__and2_4 _17516_ (.A(\cs_registers_i.mhpmcounter[1874] ),
    .B(_11951_),
    .X(_11954_));
 sky130_fd_sc_hd__o21ai_0 _17517_ (.A1(net3434),
    .A2(_11954_),
    .B1(_11899_),
    .Y(_11955_));
 sky130_fd_sc_hd__nand2_2 _17518_ (.A(\cs_registers_i.mhpmcounter[1874] ),
    .B(_11951_),
    .Y(_11956_));
 sky130_fd_sc_hd__o32ai_1 _17519_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(net3434),
    .A3(_11956_),
    .B1(_11333_),
    .B2(_11888_),
    .Y(_11957_));
 sky130_fd_sc_hd__a21o_1 _17520_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(_11955_),
    .B1(_11957_),
    .X(_00091_));
 sky130_fd_sc_hd__a21oi_1 _17521_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(net3435),
    .B1(net3490),
    .Y(_11958_));
 sky130_fd_sc_hd__nor3b_1 _17522_ (.A(_11930_),
    .B(_11958_),
    .C_N(\cs_registers_i.mhpmcounter[1857] ),
    .Y(_11959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_764 ();
 sky130_fd_sc_hd__a21oi_1 _17524_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(net3435),
    .B1(\cs_registers_i.mhpmcounter[1857] ),
    .Y(_11961_));
 sky130_fd_sc_hd__o22ai_1 _17525_ (.A1(_11354_),
    .A2(_11888_),
    .B1(_11959_),
    .B2(_11961_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_1 _17526_ (.A(\cs_registers_i.mhpmcounter[1875] ),
    .B(_11954_),
    .Y(_11962_));
 sky130_fd_sc_hd__o32a_1 _17527_ (.A1(\cs_registers_i.mhpmcounter[1876] ),
    .A2(net3434),
    .A3(_11962_),
    .B1(_11369_),
    .B2(_11888_),
    .X(_11963_));
 sky130_fd_sc_hd__a21oi_1 _17528_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(_11954_),
    .B1(net3434),
    .Y(_11964_));
 sky130_fd_sc_hd__o21ai_0 _17529_ (.A1(_11918_),
    .A2(_11964_),
    .B1(\cs_registers_i.mhpmcounter[1876] ),
    .Y(_11965_));
 sky130_fd_sc_hd__nand2_1 _17530_ (.A(_11963_),
    .B(_11965_),
    .Y(_00093_));
 sky130_fd_sc_hd__and3_4 _17531_ (.A(\cs_registers_i.mhpmcounter[1875] ),
    .B(\cs_registers_i.mhpmcounter[1876] ),
    .C(_11954_),
    .X(_11966_));
 sky130_fd_sc_hd__nand3b_1 _17532_ (.A_N(\cs_registers_i.mhpmcounter[1877] ),
    .B(net3438),
    .C(_11966_),
    .Y(_11967_));
 sky130_fd_sc_hd__nor2_1 _17533_ (.A(net3434),
    .B(_11966_),
    .Y(_11968_));
 sky130_fd_sc_hd__o21ai_0 _17534_ (.A1(_11918_),
    .A2(_11968_),
    .B1(\cs_registers_i.mhpmcounter[1877] ),
    .Y(_11969_));
 sky130_fd_sc_hd__o211ai_1 _17535_ (.A1(net3494),
    .A2(_11888_),
    .B1(_11967_),
    .C1(_11969_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand4b_1 _17536_ (.A_N(\cs_registers_i.mhpmcounter[1878] ),
    .B(net3438),
    .C(_11966_),
    .D(\cs_registers_i.mhpmcounter[1877] ),
    .Y(_11970_));
 sky130_fd_sc_hd__a21oi_1 _17537_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(_11966_),
    .B1(net3434),
    .Y(_11971_));
 sky130_fd_sc_hd__o21ai_0 _17538_ (.A1(_11918_),
    .A2(_11971_),
    .B1(\cs_registers_i.mhpmcounter[1878] ),
    .Y(_11972_));
 sky130_fd_sc_hd__o211ai_1 _17539_ (.A1(net3493),
    .A2(_11888_),
    .B1(_11970_),
    .C1(_11972_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand3_2 _17540_ (.A(\cs_registers_i.mhpmcounter[1876] ),
    .B(\cs_registers_i.mhpmcounter[1877] ),
    .C(\cs_registers_i.mhpmcounter[1878] ),
    .Y(_11973_));
 sky130_fd_sc_hd__nor2_2 _17541_ (.A(_11962_),
    .B(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__nand3b_1 _17542_ (.A_N(\cs_registers_i.mhpmcounter[1879] ),
    .B(net3438),
    .C(_11974_),
    .Y(_11975_));
 sky130_fd_sc_hd__nor2_1 _17543_ (.A(net3434),
    .B(_11974_),
    .Y(_11976_));
 sky130_fd_sc_hd__o21ai_0 _17544_ (.A1(_11918_),
    .A2(_11976_),
    .B1(\cs_registers_i.mhpmcounter[1879] ),
    .Y(_11977_));
 sky130_fd_sc_hd__o211ai_1 _17545_ (.A1(net3492),
    .A2(_11888_),
    .B1(_11975_),
    .C1(_11977_),
    .Y(_00096_));
 sky130_fd_sc_hd__nand4b_1 _17546_ (.A_N(\cs_registers_i.mhpmcounter[1880] ),
    .B(net3438),
    .C(_11974_),
    .D(\cs_registers_i.mhpmcounter[1879] ),
    .Y(_11978_));
 sky130_fd_sc_hd__a21oi_1 _17547_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_11974_),
    .B1(net3434),
    .Y(_11979_));
 sky130_fd_sc_hd__o21ai_0 _17548_ (.A1(_11918_),
    .A2(_11979_),
    .B1(\cs_registers_i.mhpmcounter[1880] ),
    .Y(_11980_));
 sky130_fd_sc_hd__o211ai_1 _17549_ (.A1(net3483),
    .A2(_11888_),
    .B1(_11978_),
    .C1(_11980_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand3_1 _17550_ (.A(\cs_registers_i.mhpmcounter[1879] ),
    .B(\cs_registers_i.mhpmcounter[1880] ),
    .C(_11974_),
    .Y(_11981_));
 sky130_fd_sc_hd__a21oi_1 _17551_ (.A1(net3438),
    .A2(_11981_),
    .B1(_11918_),
    .Y(_11982_));
 sky130_fd_sc_hd__o32a_1 _17552_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(net3434),
    .A3(_11981_),
    .B1(_11457_),
    .B2(_11888_),
    .X(_11983_));
 sky130_fd_sc_hd__o21ai_0 _17553_ (.A1(_11445_),
    .A2(_11982_),
    .B1(_11983_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand4_1 _17554_ (.A(\cs_registers_i.mhpmcounter[1875] ),
    .B(\cs_registers_i.mhpmcounter[1879] ),
    .C(\cs_registers_i.mhpmcounter[1880] ),
    .D(\cs_registers_i.mhpmcounter[1881] ),
    .Y(_11984_));
 sky130_fd_sc_hd__nor3_4 _17555_ (.A(_11956_),
    .B(_11973_),
    .C(_11984_),
    .Y(_11985_));
 sky130_fd_sc_hd__o211a_1 _17556_ (.A1(net3434),
    .A2(_11985_),
    .B1(net3428),
    .C1(\cs_registers_i.mhpmcounter[1882] ),
    .X(_11986_));
 sky130_fd_sc_hd__a21oi_1 _17557_ (.A1(net3438),
    .A2(_11985_),
    .B1(\cs_registers_i.mhpmcounter[1882] ),
    .Y(_11987_));
 sky130_fd_sc_hd__o22ai_1 _17558_ (.A1(net3482),
    .A2(_11888_),
    .B1(_11986_),
    .B2(_11987_),
    .Y(_00099_));
 sky130_fd_sc_hd__and2_4 _17559_ (.A(\cs_registers_i.mhpmcounter[1882] ),
    .B(_11985_),
    .X(_11988_));
 sky130_fd_sc_hd__o211a_1 _17560_ (.A1(net3434),
    .A2(_11988_),
    .B1(net3428),
    .C1(\cs_registers_i.mhpmcounter[1883] ),
    .X(_11989_));
 sky130_fd_sc_hd__a21oi_1 _17561_ (.A1(net3438),
    .A2(_11988_),
    .B1(\cs_registers_i.mhpmcounter[1883] ),
    .Y(_11990_));
 sky130_fd_sc_hd__o22ai_1 _17562_ (.A1(net3481),
    .A2(_11888_),
    .B1(_11989_),
    .B2(_11990_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand4b_1 _17563_ (.A_N(\cs_registers_i.mhpmcounter[1884] ),
    .B(net3438),
    .C(_11988_),
    .D(\cs_registers_i.mhpmcounter[1883] ),
    .Y(_11991_));
 sky130_fd_sc_hd__a21oi_1 _17564_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_11988_),
    .B1(net3434),
    .Y(_11992_));
 sky130_fd_sc_hd__o21ai_0 _17565_ (.A1(_11918_),
    .A2(_11992_),
    .B1(\cs_registers_i.mhpmcounter[1884] ),
    .Y(_11993_));
 sky130_fd_sc_hd__o211ai_1 _17566_ (.A1(net3480),
    .A2(_11888_),
    .B1(_11991_),
    .C1(_11993_),
    .Y(_00101_));
 sky130_fd_sc_hd__and3_4 _17567_ (.A(\cs_registers_i.mhpmcounter[1883] ),
    .B(\cs_registers_i.mhpmcounter[1884] ),
    .C(_11988_),
    .X(_11994_));
 sky130_fd_sc_hd__nand3b_1 _17568_ (.A_N(\cs_registers_i.mhpmcounter[1885] ),
    .B(net3438),
    .C(_11994_),
    .Y(_11995_));
 sky130_fd_sc_hd__nor2_1 _17569_ (.A(net3434),
    .B(_11994_),
    .Y(_11996_));
 sky130_fd_sc_hd__o21ai_0 _17570_ (.A1(_11918_),
    .A2(_11996_),
    .B1(\cs_registers_i.mhpmcounter[1885] ),
    .Y(_11997_));
 sky130_fd_sc_hd__o211ai_1 _17571_ (.A1(net3479),
    .A2(_11888_),
    .B1(_11995_),
    .C1(_11997_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand3_1 _17572_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .C(net3435),
    .Y(_11998_));
 sky130_fd_sc_hd__xnor2_1 _17573_ (.A(\cs_registers_i.mhpmcounter[1858] ),
    .B(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand2_1 _17574_ (.A(_11888_),
    .B(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__o21ai_0 _17575_ (.A1(_11082_),
    .A2(_11888_),
    .B1(_12000_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand4b_1 _17576_ (.A_N(\cs_registers_i.mhpmcounter[1886] ),
    .B(net3438),
    .C(_11994_),
    .D(\cs_registers_i.mhpmcounter[1885] ),
    .Y(_12001_));
 sky130_fd_sc_hd__a21oi_1 _17577_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(_11994_),
    .B1(net3434),
    .Y(_12002_));
 sky130_fd_sc_hd__o21ai_0 _17578_ (.A1(_11918_),
    .A2(_12002_),
    .B1(\cs_registers_i.mhpmcounter[1886] ),
    .Y(_12003_));
 sky130_fd_sc_hd__o211ai_1 _17579_ (.A1(_11550_),
    .A2(_11888_),
    .B1(_12001_),
    .C1(_12003_),
    .Y(_00104_));
 sky130_fd_sc_hd__inv_2 _17580_ (.A(_11985_),
    .Y(_12004_));
 sky130_fd_sc_hd__and3_4 _17581_ (.A(\cs_registers_i.mhpmcounter[1882] ),
    .B(\cs_registers_i.mhpmcounter[1883] ),
    .C(\cs_registers_i.mhpmcounter[1884] ),
    .X(_12005_));
 sky130_fd_sc_hd__nand3_4 _17582_ (.A(\cs_registers_i.mhpmcounter[1885] ),
    .B(\cs_registers_i.mhpmcounter[1886] ),
    .C(_12005_),
    .Y(_12006_));
 sky130_fd_sc_hd__nor2_2 _17583_ (.A(_12004_),
    .B(_12006_),
    .Y(_12007_));
 sky130_fd_sc_hd__o211a_1 _17584_ (.A1(_11897_),
    .A2(_12007_),
    .B1(_11899_),
    .C1(\cs_registers_i.mhpmcounter[1887] ),
    .X(_12008_));
 sky130_fd_sc_hd__a21oi_1 _17585_ (.A1(net3439),
    .A2(_12007_),
    .B1(\cs_registers_i.mhpmcounter[1887] ),
    .Y(_12009_));
 sky130_fd_sc_hd__o22ai_1 _17586_ (.A1(_11565_),
    .A2(_11888_),
    .B1(_12008_),
    .B2(_12009_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand4_1 _17587_ (.A(_11004_),
    .B(_10993_),
    .C(_10610_),
    .D(_11885_),
    .Y(_12010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_763 ();
 sky130_fd_sc_hd__and2_4 _17589_ (.A(\cs_registers_i.mhpmcounter[1887] ),
    .B(_12007_),
    .X(_12012_));
 sky130_fd_sc_hd__nand2_8 _17590_ (.A(_11897_),
    .B(net3500),
    .Y(_12013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_762 ();
 sky130_fd_sc_hd__o211a_1 _17592_ (.A1(net3490),
    .A2(_12012_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1888] ),
    .X(_12015_));
 sky130_fd_sc_hd__a21oi_1 _17593_ (.A1(net3439),
    .A2(_12012_),
    .B1(\cs_registers_i.mhpmcounter[1888] ),
    .Y(_12016_));
 sky130_fd_sc_hd__o22ai_1 _17594_ (.A1(_11042_),
    .A2(_12010_),
    .B1(_12015_),
    .B2(_12016_),
    .Y(_00106_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_759 ();
 sky130_fd_sc_hd__nand2_1 _17598_ (.A(\cs_registers_i.mhpmcounter[1888] ),
    .B(_12012_),
    .Y(_12020_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(_11916_),
    .B(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__and3_1 _17600_ (.A(\cs_registers_i.mhpmcounter[1889] ),
    .B(_12013_),
    .C(_12021_),
    .X(_12022_));
 sky130_fd_sc_hd__a31oi_1 _17601_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(net3439),
    .A3(_12012_),
    .B1(\cs_registers_i.mhpmcounter[1889] ),
    .Y(_12023_));
 sky130_fd_sc_hd__o22ai_1 _17602_ (.A1(_11354_),
    .A2(_12010_),
    .B1(_12022_),
    .B2(_12023_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3_4 _17603_ (.A(\cs_registers_i.mhpmcounter[1888] ),
    .B(\cs_registers_i.mhpmcounter[1889] ),
    .C(_12012_),
    .X(_12024_));
 sky130_fd_sc_hd__o211a_1 _17604_ (.A1(net3490),
    .A2(_12024_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1890] ),
    .X(_12025_));
 sky130_fd_sc_hd__a21oi_1 _17605_ (.A1(net3439),
    .A2(_12024_),
    .B1(\cs_registers_i.mhpmcounter[1890] ),
    .Y(_12026_));
 sky130_fd_sc_hd__o22ai_1 _17606_ (.A1(_11082_),
    .A2(_12010_),
    .B1(_12025_),
    .B2(_12026_),
    .Y(_00108_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_758 ();
 sky130_fd_sc_hd__nand2_1 _17608_ (.A(\cs_registers_i.mhpmcounter[1890] ),
    .B(_12024_),
    .Y(_12028_));
 sky130_fd_sc_hd__nand2_1 _17609_ (.A(_11916_),
    .B(_12028_),
    .Y(_12029_));
 sky130_fd_sc_hd__and3_1 _17610_ (.A(\cs_registers_i.mhpmcounter[1891] ),
    .B(_12013_),
    .C(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__a31oi_1 _17611_ (.A1(\cs_registers_i.mhpmcounter[1890] ),
    .A2(net3439),
    .A3(_12024_),
    .B1(\cs_registers_i.mhpmcounter[1891] ),
    .Y(_12031_));
 sky130_fd_sc_hd__o22ai_1 _17612_ (.A1(_11612_),
    .A2(_12010_),
    .B1(_12030_),
    .B2(_12031_),
    .Y(_00109_));
 sky130_fd_sc_hd__and3_4 _17613_ (.A(\cs_registers_i.mhpmcounter[1890] ),
    .B(\cs_registers_i.mhpmcounter[1891] ),
    .C(_12024_),
    .X(_12032_));
 sky130_fd_sc_hd__o211a_1 _17614_ (.A1(net3490),
    .A2(_12032_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1892] ),
    .X(_12033_));
 sky130_fd_sc_hd__a21oi_1 _17615_ (.A1(net3439),
    .A2(_12032_),
    .B1(\cs_registers_i.mhpmcounter[1892] ),
    .Y(_12034_));
 sky130_fd_sc_hd__o22ai_1 _17616_ (.A1(_11780_),
    .A2(_12010_),
    .B1(_12033_),
    .B2(_12034_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _17617_ (.A(\cs_registers_i.mhpmcounter[1892] ),
    .B(_12032_),
    .Y(_12035_));
 sky130_fd_sc_hd__nand2_1 _17618_ (.A(_11916_),
    .B(_12035_),
    .Y(_12036_));
 sky130_fd_sc_hd__and3_1 _17619_ (.A(\cs_registers_i.mhpmcounter[1893] ),
    .B(_12013_),
    .C(_12036_),
    .X(_12037_));
 sky130_fd_sc_hd__a31oi_1 _17620_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(net3439),
    .A3(_12032_),
    .B1(\cs_registers_i.mhpmcounter[1893] ),
    .Y(_12038_));
 sky130_fd_sc_hd__o22ai_1 _17621_ (.A1(_11647_),
    .A2(_12010_),
    .B1(_12037_),
    .B2(_12038_),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_1 _17622_ (.A(_12012_),
    .Y(_12039_));
 sky130_fd_sc_hd__and4_1 _17623_ (.A(\cs_registers_i.mhpmcounter[1890] ),
    .B(\cs_registers_i.mhpmcounter[1891] ),
    .C(\cs_registers_i.mhpmcounter[1892] ),
    .D(\cs_registers_i.mhpmcounter[1893] ),
    .X(_12040_));
 sky130_fd_sc_hd__nand3_2 _17624_ (.A(\cs_registers_i.mhpmcounter[1888] ),
    .B(\cs_registers_i.mhpmcounter[1889] ),
    .C(_12040_),
    .Y(_12041_));
 sky130_fd_sc_hd__nor2_1 _17625_ (.A(_12039_),
    .B(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__o211a_1 _17626_ (.A1(net3490),
    .A2(_12042_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1894] ),
    .X(_12043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_757 ();
 sky130_fd_sc_hd__a21oi_1 _17628_ (.A1(net3439),
    .A2(_12042_),
    .B1(\cs_registers_i.mhpmcounter[1894] ),
    .Y(_12045_));
 sky130_fd_sc_hd__o22ai_1 _17629_ (.A1(_11664_),
    .A2(net3500),
    .B1(_12043_),
    .B2(_12045_),
    .Y(_00112_));
 sky130_fd_sc_hd__and2_4 _17630_ (.A(\cs_registers_i.mhpmcounter[1894] ),
    .B(_12042_),
    .X(_12046_));
 sky130_fd_sc_hd__o211a_1 _17631_ (.A1(net3490),
    .A2(_12046_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1895] ),
    .X(_12047_));
 sky130_fd_sc_hd__a21oi_1 _17632_ (.A1(net3439),
    .A2(_12046_),
    .B1(\cs_registers_i.mhpmcounter[1895] ),
    .Y(_12048_));
 sky130_fd_sc_hd__o22ai_1 _17633_ (.A1(net3478),
    .A2(net3500),
    .B1(_12047_),
    .B2(_12048_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand4_1 _17634_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .C(\cs_registers_i.mhpmcounter[1858] ),
    .D(net3435),
    .Y(_12049_));
 sky130_fd_sc_hd__and3_1 _17635_ (.A(\cs_registers_i.mhpmcounter[1859] ),
    .B(_11916_),
    .C(_12049_),
    .X(_12050_));
 sky130_fd_sc_hd__a21oi_1 _17636_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(_11930_),
    .B1(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__o221ai_1 _17637_ (.A1(_11612_),
    .A2(_11888_),
    .B1(net3426),
    .B2(\cs_registers_i.mhpmcounter[1859] ),
    .C1(_12051_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _17638_ (.A(\cs_registers_i.mhpmcounter[1895] ),
    .B(_12046_),
    .Y(_12052_));
 sky130_fd_sc_hd__nand2_1 _17639_ (.A(_11916_),
    .B(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__and3_1 _17640_ (.A(\cs_registers_i.mhpmcounter[1896] ),
    .B(_12013_),
    .C(_12053_),
    .X(_12054_));
 sky130_fd_sc_hd__a31oi_1 _17641_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(net3439),
    .A3(_12046_),
    .B1(\cs_registers_i.mhpmcounter[1896] ),
    .Y(_12055_));
 sky130_fd_sc_hd__o22ai_1 _17642_ (.A1(_11707_),
    .A2(net3500),
    .B1(_12054_),
    .B2(_12055_),
    .Y(_00115_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_756 ();
 sky130_fd_sc_hd__nand3_1 _17644_ (.A(\cs_registers_i.mhpmcounter[1895] ),
    .B(\cs_registers_i.mhpmcounter[1896] ),
    .C(_12046_),
    .Y(_12057_));
 sky130_fd_sc_hd__nor2_1 _17645_ (.A(_11897_),
    .B(_12057_),
    .Y(_12058_));
 sky130_fd_sc_hd__nand2_1 _17646_ (.A(_11916_),
    .B(_12057_),
    .Y(_12059_));
 sky130_fd_sc_hd__nand3_1 _17647_ (.A(\cs_registers_i.mhpmcounter[1897] ),
    .B(_12013_),
    .C(_12059_),
    .Y(_12060_));
 sky130_fd_sc_hd__o21ai_0 _17648_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(_12058_),
    .B1(_12060_),
    .Y(_12061_));
 sky130_fd_sc_hd__o21ai_0 _17649_ (.A1(_11726_),
    .A2(net3500),
    .B1(_12061_),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_1 _17650_ (.A(\cs_registers_i.mhpmcounter[1897] ),
    .Y(_12062_));
 sky130_fd_sc_hd__nor2_1 _17651_ (.A(_12062_),
    .B(_12057_),
    .Y(_12063_));
 sky130_fd_sc_hd__o211a_1 _17652_ (.A1(net3490),
    .A2(_12063_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1898] ),
    .X(_12064_));
 sky130_fd_sc_hd__a21oi_1 _17653_ (.A1(net3439),
    .A2(_12063_),
    .B1(\cs_registers_i.mhpmcounter[1898] ),
    .Y(_12065_));
 sky130_fd_sc_hd__o22ai_1 _17654_ (.A1(_11145_),
    .A2(net3500),
    .B1(_12064_),
    .B2(_12065_),
    .Y(_00117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_755 ();
 sky130_fd_sc_hd__and2_4 _17656_ (.A(\cs_registers_i.mhpmcounter[1898] ),
    .B(_12063_),
    .X(_12067_));
 sky130_fd_sc_hd__o211a_1 _17657_ (.A1(net3490),
    .A2(_12067_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1899] ),
    .X(_12068_));
 sky130_fd_sc_hd__a21oi_1 _17658_ (.A1(net3439),
    .A2(_12067_),
    .B1(\cs_registers_i.mhpmcounter[1899] ),
    .Y(_12069_));
 sky130_fd_sc_hd__o22ai_1 _17659_ (.A1(_11177_),
    .A2(net3500),
    .B1(_12068_),
    .B2(_12069_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _17660_ (.A(\cs_registers_i.mhpmcounter[1899] ),
    .B(_12067_),
    .Y(_12070_));
 sky130_fd_sc_hd__nand2_1 _17661_ (.A(_11916_),
    .B(_12070_),
    .Y(_12071_));
 sky130_fd_sc_hd__and3_1 _17662_ (.A(\cs_registers_i.mhpmcounter[1900] ),
    .B(_12013_),
    .C(_12071_),
    .X(_12072_));
 sky130_fd_sc_hd__a31oi_1 _17663_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(net3439),
    .A3(_12067_),
    .B1(\cs_registers_i.mhpmcounter[1900] ),
    .Y(_12073_));
 sky130_fd_sc_hd__o22ai_1 _17664_ (.A1(_11197_),
    .A2(net3500),
    .B1(_12072_),
    .B2(_12073_),
    .Y(_00119_));
 sky130_fd_sc_hd__and3_4 _17665_ (.A(\cs_registers_i.mhpmcounter[1900] ),
    .B(\cs_registers_i.mhpmcounter[1899] ),
    .C(_12067_),
    .X(_12074_));
 sky130_fd_sc_hd__o211a_1 _17666_ (.A1(net3490),
    .A2(_12074_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1901] ),
    .X(_12075_));
 sky130_fd_sc_hd__a21oi_1 _17667_ (.A1(net3439),
    .A2(_12074_),
    .B1(\cs_registers_i.mhpmcounter[1901] ),
    .Y(_12076_));
 sky130_fd_sc_hd__o22ai_1 _17668_ (.A1(_11214_),
    .A2(net3500),
    .B1(_12075_),
    .B2(_12076_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(\cs_registers_i.mhpmcounter[1901] ),
    .B(_12074_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand2_1 _17670_ (.A(_11916_),
    .B(_12077_),
    .Y(_12078_));
 sky130_fd_sc_hd__and3_1 _17671_ (.A(\cs_registers_i.mhpmcounter[1902] ),
    .B(_12013_),
    .C(_12078_),
    .X(_12079_));
 sky130_fd_sc_hd__a31oi_1 _17672_ (.A1(\cs_registers_i.mhpmcounter[1901] ),
    .A2(net3439),
    .A3(_12074_),
    .B1(\cs_registers_i.mhpmcounter[1902] ),
    .Y(_12080_));
 sky130_fd_sc_hd__o22ai_1 _17673_ (.A1(_11235_),
    .A2(net3500),
    .B1(_12079_),
    .B2(_12080_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand4_1 _17674_ (.A(\cs_registers_i.mhpmcounter[1898] ),
    .B(\cs_registers_i.mhpmcounter[1901] ),
    .C(\cs_registers_i.mhpmcounter[1902] ),
    .D(\cs_registers_i.mhpmcounter[1887] ),
    .Y(_12081_));
 sky130_fd_sc_hd__nand2_1 _17675_ (.A(\cs_registers_i.mhpmcounter[1900] ),
    .B(\cs_registers_i.mhpmcounter[1899] ),
    .Y(_12082_));
 sky130_fd_sc_hd__nand4_1 _17676_ (.A(\cs_registers_i.mhpmcounter[1894] ),
    .B(\cs_registers_i.mhpmcounter[1895] ),
    .C(\cs_registers_i.mhpmcounter[1896] ),
    .D(\cs_registers_i.mhpmcounter[1897] ),
    .Y(_12083_));
 sky130_fd_sc_hd__or3_4 _17677_ (.A(_12081_),
    .B(_12082_),
    .C(_12083_),
    .X(_12084_));
 sky130_fd_sc_hd__nor4_2 _17678_ (.A(_12004_),
    .B(_12006_),
    .C(_12041_),
    .D(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__o211a_1 _17679_ (.A1(net3490),
    .A2(_12085_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1903] ),
    .X(_12086_));
 sky130_fd_sc_hd__a21oi_1 _17680_ (.A1(net3437),
    .A2(_12085_),
    .B1(\cs_registers_i.mhpmcounter[1903] ),
    .Y(_12087_));
 sky130_fd_sc_hd__o22ai_1 _17681_ (.A1(_11255_),
    .A2(net3500),
    .B1(_12086_),
    .B2(_12087_),
    .Y(_00122_));
 sky130_fd_sc_hd__and2_4 _17682_ (.A(\cs_registers_i.mhpmcounter[1903] ),
    .B(_12085_),
    .X(_12088_));
 sky130_fd_sc_hd__o211a_1 _17683_ (.A1(net3490),
    .A2(_12088_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1904] ),
    .X(_12089_));
 sky130_fd_sc_hd__a21oi_1 _17684_ (.A1(net3437),
    .A2(_12088_),
    .B1(\cs_registers_i.mhpmcounter[1904] ),
    .Y(_12090_));
 sky130_fd_sc_hd__o22ai_1 _17685_ (.A1(_11270_),
    .A2(net3500),
    .B1(_12089_),
    .B2(_12090_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _17686_ (.A(\cs_registers_i.mhpmcounter[1904] ),
    .B(_12088_),
    .Y(_12091_));
 sky130_fd_sc_hd__nand2_1 _17687_ (.A(_11916_),
    .B(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__and3_1 _17688_ (.A(\cs_registers_i.mhpmcounter[1905] ),
    .B(_12013_),
    .C(_12092_),
    .X(_12093_));
 sky130_fd_sc_hd__a31oi_1 _17689_ (.A1(\cs_registers_i.mhpmcounter[1904] ),
    .A2(net3437),
    .A3(_12088_),
    .B1(\cs_registers_i.mhpmcounter[1905] ),
    .Y(_12094_));
 sky130_fd_sc_hd__o22ai_1 _17690_ (.A1(_11294_),
    .A2(net3500),
    .B1(_12093_),
    .B2(_12094_),
    .Y(_00124_));
 sky130_fd_sc_hd__o21ai_0 _17691_ (.A1(net3434),
    .A2(_11903_),
    .B1(_11899_),
    .Y(_12095_));
 sky130_fd_sc_hd__nor3b_1 _17692_ (.A(\cs_registers_i.mhpmcounter[1860] ),
    .B(net3434),
    .C_N(_11903_),
    .Y(_12096_));
 sky130_fd_sc_hd__a221o_1 _17693_ (.A1(_11631_),
    .A2(_11917_),
    .B1(_12095_),
    .B2(\cs_registers_i.mhpmcounter[1860] ),
    .C1(_12096_),
    .X(_00125_));
 sky130_fd_sc_hd__and4_4 _17694_ (.A(\cs_registers_i.mhpmcounter[1903] ),
    .B(\cs_registers_i.mhpmcounter[1904] ),
    .C(\cs_registers_i.mhpmcounter[1905] ),
    .D(_12085_),
    .X(_12097_));
 sky130_fd_sc_hd__o211a_1 _17695_ (.A1(net3490),
    .A2(_12097_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1906] ),
    .X(_12098_));
 sky130_fd_sc_hd__a21oi_1 _17696_ (.A1(net3437),
    .A2(_12097_),
    .B1(\cs_registers_i.mhpmcounter[1906] ),
    .Y(_12099_));
 sky130_fd_sc_hd__o22ai_1 _17697_ (.A1(_11319_),
    .A2(net3500),
    .B1(_12098_),
    .B2(_12099_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _17698_ (.A(\cs_registers_i.mhpmcounter[1906] ),
    .B(_12097_),
    .Y(_12100_));
 sky130_fd_sc_hd__nand2_1 _17699_ (.A(_11916_),
    .B(_12100_),
    .Y(_12101_));
 sky130_fd_sc_hd__and3_1 _17700_ (.A(\cs_registers_i.mhpmcounter[1907] ),
    .B(_12013_),
    .C(_12101_),
    .X(_12102_));
 sky130_fd_sc_hd__a31oi_1 _17701_ (.A1(\cs_registers_i.mhpmcounter[1906] ),
    .A2(net3437),
    .A3(_12097_),
    .B1(\cs_registers_i.mhpmcounter[1907] ),
    .Y(_12103_));
 sky130_fd_sc_hd__o22ai_1 _17702_ (.A1(_11333_),
    .A2(net3500),
    .B1(_12102_),
    .B2(_12103_),
    .Y(_00127_));
 sky130_fd_sc_hd__and3_4 _17703_ (.A(\cs_registers_i.mhpmcounter[1906] ),
    .B(\cs_registers_i.mhpmcounter[1907] ),
    .C(_12097_),
    .X(_12104_));
 sky130_fd_sc_hd__o211a_1 _17704_ (.A1(net3490),
    .A2(_12104_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1908] ),
    .X(_12105_));
 sky130_fd_sc_hd__a21oi_1 _17705_ (.A1(net3438),
    .A2(_12104_),
    .B1(\cs_registers_i.mhpmcounter[1908] ),
    .Y(_12106_));
 sky130_fd_sc_hd__o22ai_1 _17706_ (.A1(_11369_),
    .A2(net3500),
    .B1(_12105_),
    .B2(_12106_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(\cs_registers_i.mhpmcounter[1908] ),
    .B(_12104_),
    .Y(_12107_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(_11916_),
    .B(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__and3_1 _17709_ (.A(\cs_registers_i.mhpmcounter[1909] ),
    .B(_12013_),
    .C(_12108_),
    .X(_12109_));
 sky130_fd_sc_hd__a31oi_1 _17710_ (.A1(\cs_registers_i.mhpmcounter[1908] ),
    .A2(net3438),
    .A3(_12104_),
    .B1(\cs_registers_i.mhpmcounter[1909] ),
    .Y(_12110_));
 sky130_fd_sc_hd__o22ai_1 _17711_ (.A1(net3494),
    .A2(net3500),
    .B1(_12109_),
    .B2(_12110_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand3_2 _17712_ (.A(\cs_registers_i.mhpmcounter[1908] ),
    .B(\cs_registers_i.mhpmcounter[1909] ),
    .C(_12104_),
    .Y(_12111_));
 sky130_fd_sc_hd__nor2_1 _17713_ (.A(net3434),
    .B(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__nand2_1 _17714_ (.A(_11916_),
    .B(_12111_),
    .Y(_12113_));
 sky130_fd_sc_hd__nand3_1 _17715_ (.A(\cs_registers_i.mhpmcounter[1910] ),
    .B(_12013_),
    .C(_12113_),
    .Y(_12114_));
 sky130_fd_sc_hd__o21ai_0 _17716_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(_12112_),
    .B1(_12114_),
    .Y(_12115_));
 sky130_fd_sc_hd__o21ai_0 _17717_ (.A1(net3493),
    .A2(net3500),
    .B1(_12115_),
    .Y(_00130_));
 sky130_fd_sc_hd__nor2_2 _17718_ (.A(_11395_),
    .B(_12111_),
    .Y(_12116_));
 sky130_fd_sc_hd__o211a_1 _17719_ (.A1(net3490),
    .A2(_12116_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1911] ),
    .X(_12117_));
 sky130_fd_sc_hd__a21oi_1 _17720_ (.A1(net3438),
    .A2(_12116_),
    .B1(\cs_registers_i.mhpmcounter[1911] ),
    .Y(_12118_));
 sky130_fd_sc_hd__o22ai_1 _17721_ (.A1(net3492),
    .A2(net3500),
    .B1(_12117_),
    .B2(_12118_),
    .Y(_00131_));
 sky130_fd_sc_hd__and2_4 _17722_ (.A(\cs_registers_i.mhpmcounter[1911] ),
    .B(_12116_),
    .X(_12119_));
 sky130_fd_sc_hd__o211a_1 _17723_ (.A1(net3490),
    .A2(_12119_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1912] ),
    .X(_12120_));
 sky130_fd_sc_hd__a21oi_1 _17724_ (.A1(net3438),
    .A2(_12119_),
    .B1(\cs_registers_i.mhpmcounter[1912] ),
    .Y(_12121_));
 sky130_fd_sc_hd__o22ai_1 _17725_ (.A1(net3483),
    .A2(net3500),
    .B1(_12120_),
    .B2(_12121_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _17726_ (.A(\cs_registers_i.mhpmcounter[1912] ),
    .B(_12119_),
    .Y(_12122_));
 sky130_fd_sc_hd__nand2_1 _17727_ (.A(_11916_),
    .B(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__and3_1 _17728_ (.A(\cs_registers_i.mhpmcounter[1913] ),
    .B(_12013_),
    .C(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__a31oi_1 _17729_ (.A1(\cs_registers_i.mhpmcounter[1912] ),
    .A2(net3438),
    .A3(_12119_),
    .B1(\cs_registers_i.mhpmcounter[1913] ),
    .Y(_12125_));
 sky130_fd_sc_hd__o22ai_1 _17730_ (.A1(_11457_),
    .A2(net3500),
    .B1(_12124_),
    .B2(_12125_),
    .Y(_00133_));
 sky130_fd_sc_hd__and3_4 _17731_ (.A(\cs_registers_i.mhpmcounter[1912] ),
    .B(\cs_registers_i.mhpmcounter[1913] ),
    .C(_12119_),
    .X(_12126_));
 sky130_fd_sc_hd__o211a_1 _17732_ (.A1(net3490),
    .A2(_12126_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1914] ),
    .X(_12127_));
 sky130_fd_sc_hd__a21oi_1 _17733_ (.A1(net3438),
    .A2(_12126_),
    .B1(\cs_registers_i.mhpmcounter[1914] ),
    .Y(_12128_));
 sky130_fd_sc_hd__o22ai_1 _17734_ (.A1(net3482),
    .A2(net3500),
    .B1(_12127_),
    .B2(_12128_),
    .Y(_00134_));
 sky130_fd_sc_hd__nand2_1 _17735_ (.A(\cs_registers_i.mhpmcounter[1914] ),
    .B(_12126_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_11916_),
    .B(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__and3_1 _17737_ (.A(\cs_registers_i.mhpmcounter[1915] ),
    .B(_12013_),
    .C(_12130_),
    .X(_12131_));
 sky130_fd_sc_hd__a31oi_1 _17738_ (.A1(\cs_registers_i.mhpmcounter[1914] ),
    .A2(net3438),
    .A3(_12126_),
    .B1(\cs_registers_i.mhpmcounter[1915] ),
    .Y(_12132_));
 sky130_fd_sc_hd__o22ai_1 _17739_ (.A1(net3481),
    .A2(net3500),
    .B1(_12131_),
    .B2(_12132_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand4b_1 _17740_ (.A_N(\cs_registers_i.mhpmcounter[1861] ),
    .B(net3438),
    .C(_11903_),
    .D(\cs_registers_i.mhpmcounter[1860] ),
    .Y(_12133_));
 sky130_fd_sc_hd__a21oi_1 _17741_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(_11903_),
    .B1(net3434),
    .Y(_12134_));
 sky130_fd_sc_hd__o21ai_0 _17742_ (.A1(_11918_),
    .A2(_12134_),
    .B1(\cs_registers_i.mhpmcounter[1861] ),
    .Y(_12135_));
 sky130_fd_sc_hd__o211ai_1 _17743_ (.A1(_11647_),
    .A2(_11888_),
    .B1(_12133_),
    .C1(_12135_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand3_2 _17744_ (.A(\cs_registers_i.mhpmcounter[1914] ),
    .B(\cs_registers_i.mhpmcounter[1915] ),
    .C(_12126_),
    .Y(_12136_));
 sky130_fd_sc_hd__nor2_1 _17745_ (.A(_11897_),
    .B(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(_11916_),
    .B(_12136_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand3_1 _17747_ (.A(\cs_registers_i.mhpmcounter[1916] ),
    .B(_12013_),
    .C(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21ai_0 _17748_ (.A1(\cs_registers_i.mhpmcounter[1916] ),
    .A2(_12137_),
    .B1(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__o21ai_0 _17749_ (.A1(net3480),
    .A2(net3500),
    .B1(_12140_),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_1 _17750_ (.A(\cs_registers_i.mhpmcounter[1916] ),
    .Y(_12141_));
 sky130_fd_sc_hd__nor2_2 _17751_ (.A(_12141_),
    .B(_12136_),
    .Y(_12142_));
 sky130_fd_sc_hd__o211a_1 _17752_ (.A1(net3490),
    .A2(_12142_),
    .B1(_12013_),
    .C1(\cs_registers_i.mhpmcounter[1917] ),
    .X(_12143_));
 sky130_fd_sc_hd__a21oi_1 _17753_ (.A1(net3437),
    .A2(_12142_),
    .B1(\cs_registers_i.mhpmcounter[1917] ),
    .Y(_12144_));
 sky130_fd_sc_hd__o22ai_1 _17754_ (.A1(net3479),
    .A2(net3500),
    .B1(_12143_),
    .B2(_12144_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(\cs_registers_i.mhpmcounter[1917] ),
    .B(_12142_),
    .Y(_12145_));
 sky130_fd_sc_hd__nand2_1 _17756_ (.A(_11916_),
    .B(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__and3_1 _17757_ (.A(\cs_registers_i.mhpmcounter[1918] ),
    .B(_12013_),
    .C(_12146_),
    .X(_12147_));
 sky130_fd_sc_hd__a31oi_1 _17758_ (.A1(\cs_registers_i.mhpmcounter[1917] ),
    .A2(net3437),
    .A3(_12142_),
    .B1(\cs_registers_i.mhpmcounter[1918] ),
    .Y(_12148_));
 sky130_fd_sc_hd__o22ai_1 _17759_ (.A1(_11550_),
    .A2(net3500),
    .B1(_12147_),
    .B2(_12148_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand3_1 _17760_ (.A(\cs_registers_i.mhpmcounter[1917] ),
    .B(\cs_registers_i.mhpmcounter[1918] ),
    .C(_12142_),
    .Y(_12149_));
 sky130_fd_sc_hd__nand2_1 _17761_ (.A(_11916_),
    .B(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__and3_1 _17762_ (.A(\cs_registers_i.mhpmcounter[1919] ),
    .B(_12013_),
    .C(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__a41oi_1 _17763_ (.A1(\cs_registers_i.mhpmcounter[1917] ),
    .A2(\cs_registers_i.mhpmcounter[1918] ),
    .A3(net3437),
    .A4(_12142_),
    .B1(\cs_registers_i.mhpmcounter[1919] ),
    .Y(_12152_));
 sky130_fd_sc_hd__o22ai_1 _17764_ (.A1(_11565_),
    .A2(net3500),
    .B1(_12151_),
    .B2(_12152_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(net3435),
    .B(_11904_),
    .Y(_12153_));
 sky130_fd_sc_hd__and3_1 _17766_ (.A(\cs_registers_i.mhpmcounter[1862] ),
    .B(_11916_),
    .C(_12153_),
    .X(_12154_));
 sky130_fd_sc_hd__a21oi_1 _17767_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_11930_),
    .B1(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__o221ai_1 _17768_ (.A1(_11664_),
    .A2(_11888_),
    .B1(_12153_),
    .B2(\cs_registers_i.mhpmcounter[1862] ),
    .C1(_12155_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand3b_1 _17769_ (.A_N(\cs_registers_i.mhpmcounter[1863] ),
    .B(net3435),
    .C(_11911_),
    .Y(_12156_));
 sky130_fd_sc_hd__nor2_1 _17770_ (.A(_11897_),
    .B(_11911_),
    .Y(_12157_));
 sky130_fd_sc_hd__o21ai_0 _17771_ (.A1(_11918_),
    .A2(_12157_),
    .B1(\cs_registers_i.mhpmcounter[1863] ),
    .Y(_12158_));
 sky130_fd_sc_hd__o211ai_1 _17772_ (.A1(net3478),
    .A2(_11888_),
    .B1(_12156_),
    .C1(_12158_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _17773_ (.A(net3435),
    .B(_11905_),
    .Y(_12159_));
 sky130_fd_sc_hd__and3_1 _17774_ (.A(\cs_registers_i.mhpmcounter[1864] ),
    .B(_11916_),
    .C(_12159_),
    .X(_12160_));
 sky130_fd_sc_hd__a21oi_1 _17775_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_11930_),
    .B1(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__o221ai_1 _17776_ (.A1(_11707_),
    .A2(_11888_),
    .B1(_12159_),
    .B2(\cs_registers_i.mhpmcounter[1864] ),
    .C1(_12161_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _17777_ (.A(\cs_registers_i.mhpmcounter[1864] ),
    .B(_11905_),
    .Y(_12162_));
 sky130_fd_sc_hd__and3_1 _17778_ (.A(\cs_registers_i.mhpmcounter[1865] ),
    .B(net3436),
    .C(_12162_),
    .X(_12163_));
 sky130_fd_sc_hd__nor3_1 _17779_ (.A(\cs_registers_i.mhpmcounter[1865] ),
    .B(net3434),
    .C(_12162_),
    .Y(_12164_));
 sky130_fd_sc_hd__a211oi_1 _17780_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_11918_),
    .B1(_12163_),
    .C1(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__o21ai_0 _17781_ (.A1(_11726_),
    .A2(_11888_),
    .B1(_12165_),
    .Y(_00144_));
 sky130_fd_sc_hd__nor2_2 _17782_ (.A(_10500_),
    .B(_10784_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand2_4 _17783_ (.A(_10796_),
    .B(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_2 _17784_ (.A(_10783_),
    .B(_10784_),
    .Y(_12168_));
 sky130_fd_sc_hd__inv_2 _17785_ (.A(_10823_),
    .Y(_12169_));
 sky130_fd_sc_hd__nor3_4 _17786_ (.A(_10495_),
    .B(_10782_),
    .C(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__nand2_8 _17787_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(_10798_),
    .Y(_12171_));
 sky130_fd_sc_hd__nor2_4 _17788_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__o21ai_4 _17789_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(net60),
    .B1(_12172_),
    .Y(_12173_));
 sky130_fd_sc_hd__nor2b_4 _17790_ (.A(net3573),
    .B_N(_12173_),
    .Y(_12174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_754 ();
 sky130_fd_sc_hd__and2_4 _17792_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(_10798_),
    .X(_12176_));
 sky130_fd_sc_hd__nand4_1 _17793_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10501_),
    .C(_10791_),
    .D(_12176_),
    .Y(_12177_));
 sky130_fd_sc_hd__o211ai_1 _17794_ (.A1(_10793_),
    .A2(_12168_),
    .B1(_12174_),
    .C1(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__nor2_1 _17795_ (.A(net3950),
    .B(net3545),
    .Y(_12179_));
 sky130_fd_sc_hd__o21ai_2 _17796_ (.A1(_10503_),
    .A2(_10512_),
    .B1(_12166_),
    .Y(_12180_));
 sky130_fd_sc_hd__nor3_4 _17797_ (.A(_10505_),
    .B(_10508_),
    .C(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_751 ();
 sky130_fd_sc_hd__a221oi_1 _17801_ (.A1(\cs_registers_i.mstatus_q[2] ),
    .A2(_10642_),
    .B1(_12181_),
    .B2(\cs_registers_i.dcsr_q[0] ),
    .C1(_12167_),
    .Y(_12185_));
 sky130_fd_sc_hd__a21oi_1 _17802_ (.A1(_12167_),
    .A2(_12179_),
    .B1(_12185_),
    .Y(_00145_));
 sky130_fd_sc_hd__nor2_1 _17803_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(net3545),
    .Y(_12186_));
 sky130_fd_sc_hd__a221oi_1 _17804_ (.A1(\cs_registers_i.mstatus_q[3] ),
    .A2(_10642_),
    .B1(_12181_),
    .B2(\cs_registers_i.dcsr_q[1] ),
    .C1(_12167_),
    .Y(_12187_));
 sky130_fd_sc_hd__a21oi_1 _17805_ (.A1(_12167_),
    .A2(_12186_),
    .B1(_12187_),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_8 _17806_ (.A(_12177_),
    .B(_12173_),
    .Y(_12188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_750 ();
 sky130_fd_sc_hd__a21oi_1 _17808_ (.A1(_11885_),
    .A2(_11030_),
    .B1(\cs_registers_i.dcsr_q[0] ),
    .Y(_12190_));
 sky130_fd_sc_hd__nand2_8 _17809_ (.A(net3501),
    .B(_11342_),
    .Y(_12191_));
 sky130_fd_sc_hd__and3b_4 _17810_ (.A_N(_12191_),
    .B(_11042_),
    .C(_11354_),
    .X(_12192_));
 sky130_fd_sc_hd__nand2_1 _17811_ (.A(net3950),
    .B(_12188_),
    .Y(_12193_));
 sky130_fd_sc_hd__o31ai_1 _17812_ (.A1(_12188_),
    .A2(_12190_),
    .A3(_12192_),
    .B1(_12193_),
    .Y(_00147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_749 ();
 sky130_fd_sc_hd__nand2_1 _17814_ (.A(\cs_registers_i.dcsr_q[11] ),
    .B(_12191_),
    .Y(_12195_));
 sky130_fd_sc_hd__o21ai_0 _17815_ (.A1(_11177_),
    .A2(_12191_),
    .B1(_12195_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _17816_ (.A(\cs_registers_i.dcsr_q[12] ),
    .B(_12191_),
    .Y(_12196_));
 sky130_fd_sc_hd__o21ai_0 _17817_ (.A1(_11197_),
    .A2(_12191_),
    .B1(_12196_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand2_1 _17818_ (.A(\cs_registers_i.dcsr_q[13] ),
    .B(_12191_),
    .Y(_12197_));
 sky130_fd_sc_hd__o21ai_0 _17819_ (.A1(_11214_),
    .A2(_12191_),
    .B1(_12197_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2_1 _17820_ (.A(\cs_registers_i.dcsr_q[15] ),
    .B(_12191_),
    .Y(_12198_));
 sky130_fd_sc_hd__o21ai_0 _17821_ (.A1(_11255_),
    .A2(_12191_),
    .B1(_12198_),
    .Y(_00151_));
 sky130_fd_sc_hd__a21oi_1 _17822_ (.A1(_11885_),
    .A2(_11030_),
    .B1(\cs_registers_i.dcsr_q[1] ),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_1 _17823_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(_12188_),
    .Y(_12200_));
 sky130_fd_sc_hd__o31ai_1 _17824_ (.A1(_12188_),
    .A2(_12192_),
    .A3(_12199_),
    .B1(_12200_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _17825_ (.A(\cs_registers_i.dcsr_q[2] ),
    .B(_12191_),
    .Y(_12201_));
 sky130_fd_sc_hd__o21ai_0 _17826_ (.A1(_11082_),
    .A2(_12191_),
    .B1(_12201_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2_1 _17827_ (.A(\cs_registers_i.dcsr_q[6] ),
    .B(_12188_),
    .Y(_12202_));
 sky130_fd_sc_hd__a21oi_1 _17828_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_12172_),
    .B1(_12202_),
    .Y(_00154_));
 sky130_fd_sc_hd__a22oi_1 _17829_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_12177_),
    .B1(_12172_),
    .B2(net60),
    .Y(_12203_));
 sky130_fd_sc_hd__a21oi_1 _17830_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_12172_),
    .B1(_12203_),
    .Y(_00155_));
 sky130_fd_sc_hd__a32o_1 _17831_ (.A1(\cs_registers_i.dcsr_q[8] ),
    .A2(_12177_),
    .A3(_12173_),
    .B1(_12172_),
    .B2(\cs_registers_i.dcsr_q[2] ),
    .X(_00156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_746 ();
 sky130_fd_sc_hd__mux2i_1 _17835_ (.A0(\cs_registers_i.pc_if_i[10] ),
    .A1(\cs_registers_i.pc_id_i[10] ),
    .S(_12174_),
    .Y(_12207_));
 sky130_fd_sc_hd__nand2_8 _17836_ (.A(net3501),
    .B(_11221_),
    .Y(_12208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_744 ();
 sky130_fd_sc_hd__nor2_1 _17839_ (.A(_11145_),
    .B(_12208_),
    .Y(_12211_));
 sky130_fd_sc_hd__a211oi_1 _17840_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(_12208_),
    .B1(_12211_),
    .C1(_12188_),
    .Y(_12212_));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_12188_),
    .A2(_12207_),
    .B1(_12212_),
    .Y(_00157_));
 sky130_fd_sc_hd__mux2i_2 _17842_ (.A0(\cs_registers_i.pc_if_i[11] ),
    .A1(\cs_registers_i.pc_id_i[11] ),
    .S(_12174_),
    .Y(_12213_));
 sky130_fd_sc_hd__nor2_1 _17843_ (.A(_11177_),
    .B(_12208_),
    .Y(_12214_));
 sky130_fd_sc_hd__a211oi_1 _17844_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_12208_),
    .B1(_12214_),
    .C1(_12188_),
    .Y(_12215_));
 sky130_fd_sc_hd__a21oi_1 _17845_ (.A1(_12188_),
    .A2(_12213_),
    .B1(_12215_),
    .Y(_00158_));
 sky130_fd_sc_hd__mux2i_1 _17846_ (.A0(\cs_registers_i.pc_if_i[12] ),
    .A1(\cs_registers_i.pc_id_i[12] ),
    .S(_12174_),
    .Y(_12216_));
 sky130_fd_sc_hd__nor2_1 _17847_ (.A(_11197_),
    .B(_12208_),
    .Y(_12217_));
 sky130_fd_sc_hd__a211oi_1 _17848_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_12208_),
    .B1(_12217_),
    .C1(_12188_),
    .Y(_12218_));
 sky130_fd_sc_hd__a21oi_1 _17849_ (.A1(_12188_),
    .A2(_12216_),
    .B1(_12218_),
    .Y(_00159_));
 sky130_fd_sc_hd__mux2i_1 _17850_ (.A0(\cs_registers_i.pc_if_i[13] ),
    .A1(\cs_registers_i.pc_id_i[13] ),
    .S(net3564),
    .Y(_12219_));
 sky130_fd_sc_hd__nor2_1 _17851_ (.A(_11214_),
    .B(_12208_),
    .Y(_12220_));
 sky130_fd_sc_hd__a211oi_1 _17852_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_12208_),
    .B1(_12220_),
    .C1(_12188_),
    .Y(_12221_));
 sky130_fd_sc_hd__a21oi_1 _17853_ (.A1(_12188_),
    .A2(_12219_),
    .B1(_12221_),
    .Y(_00160_));
 sky130_fd_sc_hd__mux2i_2 _17854_ (.A0(\cs_registers_i.pc_if_i[14] ),
    .A1(\cs_registers_i.pc_id_i[14] ),
    .S(_12174_),
    .Y(_12222_));
 sky130_fd_sc_hd__nor2_1 _17855_ (.A(_11235_),
    .B(_12208_),
    .Y(_12223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_743 ();
 sky130_fd_sc_hd__a211oi_1 _17857_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_12208_),
    .B1(_12223_),
    .C1(_12188_),
    .Y(_12225_));
 sky130_fd_sc_hd__a21oi_1 _17858_ (.A1(_12188_),
    .A2(_12222_),
    .B1(_12225_),
    .Y(_00161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_742 ();
 sky130_fd_sc_hd__mux2i_1 _17860_ (.A0(\cs_registers_i.pc_if_i[15] ),
    .A1(\cs_registers_i.pc_id_i[15] ),
    .S(net3563),
    .Y(_12227_));
 sky130_fd_sc_hd__nor2_1 _17861_ (.A(_11255_),
    .B(_12208_),
    .Y(_12228_));
 sky130_fd_sc_hd__a211oi_1 _17862_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_12208_),
    .B1(_12228_),
    .C1(_12188_),
    .Y(_12229_));
 sky130_fd_sc_hd__a21oi_1 _17863_ (.A1(_12188_),
    .A2(_12227_),
    .B1(_12229_),
    .Y(_00162_));
 sky130_fd_sc_hd__mux2i_1 _17864_ (.A0(\cs_registers_i.pc_if_i[16] ),
    .A1(\cs_registers_i.pc_id_i[16] ),
    .S(net3564),
    .Y(_12230_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_11270_),
    .B(_12208_),
    .Y(_12231_));
 sky130_fd_sc_hd__a211oi_1 _17866_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(_12208_),
    .B1(_12231_),
    .C1(_12188_),
    .Y(_12232_));
 sky130_fd_sc_hd__a21oi_1 _17867_ (.A1(_12188_),
    .A2(_12230_),
    .B1(_12232_),
    .Y(_00163_));
 sky130_fd_sc_hd__mux2i_1 _17868_ (.A0(\cs_registers_i.pc_if_i[17] ),
    .A1(\cs_registers_i.pc_id_i[17] ),
    .S(net3564),
    .Y(_12233_));
 sky130_fd_sc_hd__nor2_1 _17869_ (.A(_11294_),
    .B(_12208_),
    .Y(_12234_));
 sky130_fd_sc_hd__a211oi_1 _17870_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_12208_),
    .B1(_12234_),
    .C1(_12188_),
    .Y(_12235_));
 sky130_fd_sc_hd__a21oi_1 _17871_ (.A1(_12188_),
    .A2(_12233_),
    .B1(_12235_),
    .Y(_00164_));
 sky130_fd_sc_hd__mux2i_4 _17872_ (.A0(\cs_registers_i.pc_if_i[18] ),
    .A1(\cs_registers_i.pc_id_i[18] ),
    .S(net3564),
    .Y(_12236_));
 sky130_fd_sc_hd__nor2_1 _17873_ (.A(_11319_),
    .B(_12208_),
    .Y(_12237_));
 sky130_fd_sc_hd__a211oi_1 _17874_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(_12208_),
    .B1(_12237_),
    .C1(_12188_),
    .Y(_12238_));
 sky130_fd_sc_hd__a21oi_1 _17875_ (.A1(_12188_),
    .A2(_12236_),
    .B1(_12238_),
    .Y(_00165_));
 sky130_fd_sc_hd__mux2i_4 _17876_ (.A0(\cs_registers_i.pc_if_i[19] ),
    .A1(\cs_registers_i.pc_id_i[19] ),
    .S(net3564),
    .Y(_12239_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_741 ();
 sky130_fd_sc_hd__nor2_1 _17878_ (.A(_11333_),
    .B(_12208_),
    .Y(_12241_));
 sky130_fd_sc_hd__a211oi_1 _17879_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_12208_),
    .B1(_12241_),
    .C1(_12188_),
    .Y(_12242_));
 sky130_fd_sc_hd__a21oi_1 _17880_ (.A1(_12188_),
    .A2(_12239_),
    .B1(_12242_),
    .Y(_00166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_738 ();
 sky130_fd_sc_hd__mux2i_1 _17884_ (.A0(net3948),
    .A1(\cs_registers_i.pc_id_i[1] ),
    .S(net3564),
    .Y(_12246_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_737 ();
 sky130_fd_sc_hd__nor2_1 _17886_ (.A(_11354_),
    .B(_12208_),
    .Y(_12248_));
 sky130_fd_sc_hd__a211oi_1 _17887_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(_12208_),
    .B1(_12248_),
    .C1(_12188_),
    .Y(_12249_));
 sky130_fd_sc_hd__a21oi_1 _17888_ (.A1(_12188_),
    .A2(_12246_),
    .B1(_12249_),
    .Y(_00167_));
 sky130_fd_sc_hd__mux2i_4 _17889_ (.A0(\cs_registers_i.pc_if_i[20] ),
    .A1(\cs_registers_i.pc_id_i[20] ),
    .S(net3564),
    .Y(_12250_));
 sky130_fd_sc_hd__nor2_1 _17890_ (.A(_11369_),
    .B(_12208_),
    .Y(_12251_));
 sky130_fd_sc_hd__a211oi_1 _17891_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(_12208_),
    .B1(_12251_),
    .C1(_12188_),
    .Y(_12252_));
 sky130_fd_sc_hd__a21oi_1 _17892_ (.A1(_12188_),
    .A2(_12250_),
    .B1(_12252_),
    .Y(_00168_));
 sky130_fd_sc_hd__mux2i_1 _17893_ (.A0(\cs_registers_i.pc_if_i[21] ),
    .A1(\cs_registers_i.pc_id_i[21] ),
    .S(net3563),
    .Y(_12253_));
 sky130_fd_sc_hd__nor2_1 _17894_ (.A(_11390_),
    .B(_12208_),
    .Y(_12254_));
 sky130_fd_sc_hd__a211oi_1 _17895_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_12208_),
    .B1(_12254_),
    .C1(_12188_),
    .Y(_12255_));
 sky130_fd_sc_hd__a21oi_1 _17896_ (.A1(_12188_),
    .A2(_12253_),
    .B1(_12255_),
    .Y(_00169_));
 sky130_fd_sc_hd__mux2i_2 _17897_ (.A0(\cs_registers_i.pc_if_i[22] ),
    .A1(\cs_registers_i.pc_id_i[22] ),
    .S(net3564),
    .Y(_12256_));
 sky130_fd_sc_hd__nor2_1 _17898_ (.A(_11406_),
    .B(_12208_),
    .Y(_12257_));
 sky130_fd_sc_hd__a211oi_1 _17899_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(_12208_),
    .B1(_12257_),
    .C1(_12188_),
    .Y(_12258_));
 sky130_fd_sc_hd__a21oi_1 _17900_ (.A1(_12188_),
    .A2(_12256_),
    .B1(_12258_),
    .Y(_00170_));
 sky130_fd_sc_hd__mux2i_4 _17901_ (.A0(\cs_registers_i.pc_if_i[23] ),
    .A1(\cs_registers_i.pc_id_i[23] ),
    .S(net3564),
    .Y(_12259_));
 sky130_fd_sc_hd__nor2_1 _17902_ (.A(_11426_),
    .B(_12208_),
    .Y(_12260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_736 ();
 sky130_fd_sc_hd__a211oi_1 _17904_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_12208_),
    .B1(_12260_),
    .C1(_12188_),
    .Y(_12262_));
 sky130_fd_sc_hd__a21oi_1 _17905_ (.A1(_12188_),
    .A2(_12259_),
    .B1(_12262_),
    .Y(_00171_));
 sky130_fd_sc_hd__mux2i_1 _17906_ (.A0(\cs_registers_i.pc_if_i[24] ),
    .A1(\cs_registers_i.pc_id_i[24] ),
    .S(net3563),
    .Y(_12263_));
 sky130_fd_sc_hd__nor2_1 _17907_ (.A(_11441_),
    .B(_12208_),
    .Y(_12264_));
 sky130_fd_sc_hd__a211oi_1 _17908_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_12208_),
    .B1(_12264_),
    .C1(_12188_),
    .Y(_12265_));
 sky130_fd_sc_hd__a21oi_1 _17909_ (.A1(_12188_),
    .A2(_12263_),
    .B1(_12265_),
    .Y(_00172_));
 sky130_fd_sc_hd__mux2i_2 _17910_ (.A0(\cs_registers_i.pc_if_i[25] ),
    .A1(\cs_registers_i.pc_id_i[25] ),
    .S(net3564),
    .Y(_12266_));
 sky130_fd_sc_hd__nor2_1 _17911_ (.A(_11457_),
    .B(_12208_),
    .Y(_12267_));
 sky130_fd_sc_hd__a211oi_1 _17912_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_12208_),
    .B1(_12267_),
    .C1(_12188_),
    .Y(_12268_));
 sky130_fd_sc_hd__a21oi_1 _17913_ (.A1(_12188_),
    .A2(_12266_),
    .B1(_12268_),
    .Y(_00173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_735 ();
 sky130_fd_sc_hd__mux2i_2 _17915_ (.A0(\cs_registers_i.pc_if_i[26] ),
    .A1(net3826),
    .S(net3563),
    .Y(_12270_));
 sky130_fd_sc_hd__nor2_1 _17916_ (.A(_11476_),
    .B(_12208_),
    .Y(_12271_));
 sky130_fd_sc_hd__a211oi_1 _17917_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_12208_),
    .B1(_12271_),
    .C1(_12188_),
    .Y(_12272_));
 sky130_fd_sc_hd__a21oi_1 _17918_ (.A1(_12188_),
    .A2(_12270_),
    .B1(_12272_),
    .Y(_00174_));
 sky130_fd_sc_hd__mux2i_2 _17919_ (.A0(\cs_registers_i.pc_if_i[27] ),
    .A1(net3825),
    .S(net3563),
    .Y(_12273_));
 sky130_fd_sc_hd__nor2_1 _17920_ (.A(_11490_),
    .B(_12208_),
    .Y(_12274_));
 sky130_fd_sc_hd__a211oi_1 _17921_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_12208_),
    .B1(_12274_),
    .C1(_12188_),
    .Y(_12275_));
 sky130_fd_sc_hd__a21oi_1 _17922_ (.A1(_12188_),
    .A2(_12273_),
    .B1(_12275_),
    .Y(_00175_));
 sky130_fd_sc_hd__mux2i_2 _17923_ (.A0(\cs_registers_i.pc_if_i[28] ),
    .A1(net3824),
    .S(net3563),
    .Y(_12276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_734 ();
 sky130_fd_sc_hd__nor2_1 _17925_ (.A(_11506_),
    .B(_12208_),
    .Y(_12278_));
 sky130_fd_sc_hd__a211oi_1 _17926_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_12208_),
    .B1(_12278_),
    .C1(_12188_),
    .Y(_12279_));
 sky130_fd_sc_hd__a21oi_1 _17927_ (.A1(_12188_),
    .A2(_12276_),
    .B1(_12279_),
    .Y(_00176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_733 ();
 sky130_fd_sc_hd__mux2i_2 _17929_ (.A0(\cs_registers_i.pc_if_i[29] ),
    .A1(\cs_registers_i.pc_id_i[29] ),
    .S(net3563),
    .Y(_12281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_732 ();
 sky130_fd_sc_hd__nor2_1 _17931_ (.A(_11530_),
    .B(_12208_),
    .Y(_12283_));
 sky130_fd_sc_hd__a211oi_1 _17932_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_12208_),
    .B1(_12283_),
    .C1(_12188_),
    .Y(_12284_));
 sky130_fd_sc_hd__a21oi_1 _17933_ (.A1(_12188_),
    .A2(_12281_),
    .B1(_12284_),
    .Y(_00177_));
 sky130_fd_sc_hd__mux2i_2 _17934_ (.A0(\cs_registers_i.pc_if_i[2] ),
    .A1(\cs_registers_i.pc_id_i[2] ),
    .S(_12174_),
    .Y(_12285_));
 sky130_fd_sc_hd__nor2_1 _17935_ (.A(_11082_),
    .B(_12208_),
    .Y(_12286_));
 sky130_fd_sc_hd__a211oi_1 _17936_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_12208_),
    .B1(_12286_),
    .C1(_12188_),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_1 _17937_ (.A1(_12188_),
    .A2(_12285_),
    .B1(_12287_),
    .Y(_00178_));
 sky130_fd_sc_hd__mux2i_2 _17938_ (.A0(\cs_registers_i.pc_if_i[30] ),
    .A1(\cs_registers_i.pc_id_i[30] ),
    .S(net3564),
    .Y(_12288_));
 sky130_fd_sc_hd__nor2_1 _17939_ (.A(_11550_),
    .B(_12208_),
    .Y(_12289_));
 sky130_fd_sc_hd__a211oi_1 _17940_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(_12208_),
    .B1(_12289_),
    .C1(_12188_),
    .Y(_12290_));
 sky130_fd_sc_hd__a21oi_1 _17941_ (.A1(_12188_),
    .A2(_12288_),
    .B1(_12290_),
    .Y(_00179_));
 sky130_fd_sc_hd__mux2i_1 _17942_ (.A0(\cs_registers_i.pc_if_i[31] ),
    .A1(\cs_registers_i.pc_id_i[31] ),
    .S(net3564),
    .Y(_12291_));
 sky130_fd_sc_hd__nor2_1 _17943_ (.A(_11565_),
    .B(_12208_),
    .Y(_12292_));
 sky130_fd_sc_hd__a211oi_1 _17944_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_12208_),
    .B1(_12292_),
    .C1(_12188_),
    .Y(_12293_));
 sky130_fd_sc_hd__a21oi_1 _17945_ (.A1(_12188_),
    .A2(_12291_),
    .B1(_12293_),
    .Y(_00180_));
 sky130_fd_sc_hd__mux2i_4 _17946_ (.A0(\cs_registers_i.pc_if_i[3] ),
    .A1(\cs_registers_i.pc_id_i[3] ),
    .S(_12174_),
    .Y(_12294_));
 sky130_fd_sc_hd__nor2_1 _17947_ (.A(_11612_),
    .B(_12208_),
    .Y(_12295_));
 sky130_fd_sc_hd__a211oi_1 _17948_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(_12208_),
    .B1(_12295_),
    .C1(_12188_),
    .Y(_12296_));
 sky130_fd_sc_hd__a21oi_1 _17949_ (.A1(_12188_),
    .A2(_12294_),
    .B1(_12296_),
    .Y(_00181_));
 sky130_fd_sc_hd__mux2i_1 _17950_ (.A0(\cs_registers_i.pc_if_i[4] ),
    .A1(\cs_registers_i.pc_id_i[4] ),
    .S(net3564),
    .Y(_12297_));
 sky130_fd_sc_hd__nor2_1 _17951_ (.A(_11780_),
    .B(_12208_),
    .Y(_12298_));
 sky130_fd_sc_hd__a211oi_1 _17952_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(_12208_),
    .B1(_12298_),
    .C1(_12188_),
    .Y(_12299_));
 sky130_fd_sc_hd__a21oi_1 _17953_ (.A1(_12188_),
    .A2(_12297_),
    .B1(_12299_),
    .Y(_00182_));
 sky130_fd_sc_hd__mux2i_2 _17954_ (.A0(\cs_registers_i.pc_if_i[5] ),
    .A1(\cs_registers_i.pc_id_i[5] ),
    .S(net3564),
    .Y(_12300_));
 sky130_fd_sc_hd__nor2_1 _17955_ (.A(_11647_),
    .B(_12208_),
    .Y(_12301_));
 sky130_fd_sc_hd__a211oi_1 _17956_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(_12208_),
    .B1(_12301_),
    .C1(_12188_),
    .Y(_12302_));
 sky130_fd_sc_hd__a21oi_1 _17957_ (.A1(_12188_),
    .A2(_12300_),
    .B1(_12302_),
    .Y(_00183_));
 sky130_fd_sc_hd__mux2i_1 _17958_ (.A0(\cs_registers_i.pc_if_i[6] ),
    .A1(\cs_registers_i.pc_id_i[6] ),
    .S(net3564),
    .Y(_12303_));
 sky130_fd_sc_hd__nor2_1 _17959_ (.A(_11664_),
    .B(_12208_),
    .Y(_12304_));
 sky130_fd_sc_hd__a211oi_1 _17960_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(_12208_),
    .B1(_12304_),
    .C1(_12188_),
    .Y(_12305_));
 sky130_fd_sc_hd__a21oi_1 _17961_ (.A1(_12188_),
    .A2(_12303_),
    .B1(_12305_),
    .Y(_00184_));
 sky130_fd_sc_hd__mux2i_1 _17962_ (.A0(\cs_registers_i.pc_if_i[7] ),
    .A1(\cs_registers_i.pc_id_i[7] ),
    .S(_12174_),
    .Y(_12306_));
 sky130_fd_sc_hd__nor2_1 _17963_ (.A(_11685_),
    .B(_12208_),
    .Y(_12307_));
 sky130_fd_sc_hd__a211oi_1 _17964_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_12208_),
    .B1(_12307_),
    .C1(_12188_),
    .Y(_12308_));
 sky130_fd_sc_hd__a21oi_1 _17965_ (.A1(_12188_),
    .A2(_12306_),
    .B1(_12308_),
    .Y(_00185_));
 sky130_fd_sc_hd__mux2i_2 _17966_ (.A0(\cs_registers_i.pc_if_i[8] ),
    .A1(net3823),
    .S(_12174_),
    .Y(_12309_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(_11707_),
    .B(_12208_),
    .Y(_12310_));
 sky130_fd_sc_hd__a211oi_1 _17968_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(_12208_),
    .B1(_12310_),
    .C1(_12188_),
    .Y(_12311_));
 sky130_fd_sc_hd__a21oi_1 _17969_ (.A1(_12188_),
    .A2(_12309_),
    .B1(_12311_),
    .Y(_00186_));
 sky130_fd_sc_hd__mux2i_2 _17970_ (.A0(\cs_registers_i.pc_if_i[9] ),
    .A1(\cs_registers_i.pc_id_i[9] ),
    .S(_12174_),
    .Y(_12312_));
 sky130_fd_sc_hd__nor2_1 _17971_ (.A(_11726_),
    .B(_12208_),
    .Y(_12313_));
 sky130_fd_sc_hd__a211oi_1 _17972_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(_12208_),
    .B1(_12313_),
    .C1(_12188_),
    .Y(_12314_));
 sky130_fd_sc_hd__a21oi_1 _17973_ (.A1(_12188_),
    .A2(_12312_),
    .B1(_12314_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_8 _17974_ (.A(net3501),
    .B(_11228_),
    .Y(_12315_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_730 ();
 sky130_fd_sc_hd__nand2_1 _17977_ (.A(\cs_registers_i.dscratch0_q[0] ),
    .B(_12315_),
    .Y(_12318_));
 sky130_fd_sc_hd__o21ai_0 _17978_ (.A1(_11042_),
    .A2(_12315_),
    .B1(_12318_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _17979_ (.A(\cs_registers_i.dscratch0_q[10] ),
    .B(_12315_),
    .Y(_12319_));
 sky130_fd_sc_hd__o21ai_0 _17980_ (.A1(_11145_),
    .A2(_12315_),
    .B1(_12319_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _17981_ (.A(\cs_registers_i.dscratch0_q[11] ),
    .B(_12315_),
    .Y(_12320_));
 sky130_fd_sc_hd__o21ai_0 _17982_ (.A1(_11177_),
    .A2(_12315_),
    .B1(_12320_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _17983_ (.A(\cs_registers_i.dscratch0_q[12] ),
    .B(_12315_),
    .Y(_12321_));
 sky130_fd_sc_hd__o21ai_0 _17984_ (.A1(_11197_),
    .A2(_12315_),
    .B1(_12321_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(\cs_registers_i.dscratch0_q[13] ),
    .B(_12315_),
    .Y(_12322_));
 sky130_fd_sc_hd__o21ai_0 _17986_ (.A1(_11214_),
    .A2(_12315_),
    .B1(_12322_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _17987_ (.A(\cs_registers_i.dscratch0_q[14] ),
    .B(_12315_),
    .Y(_12323_));
 sky130_fd_sc_hd__o21ai_0 _17988_ (.A1(_11235_),
    .A2(_12315_),
    .B1(_12323_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _17989_ (.A(\cs_registers_i.dscratch0_q[15] ),
    .B(_12315_),
    .Y(_12324_));
 sky130_fd_sc_hd__o21ai_0 _17990_ (.A1(_11255_),
    .A2(_12315_),
    .B1(_12324_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(\cs_registers_i.dscratch0_q[16] ),
    .B(_12315_),
    .Y(_12325_));
 sky130_fd_sc_hd__o21ai_0 _17992_ (.A1(_11270_),
    .A2(_12315_),
    .B1(_12325_),
    .Y(_00195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_729 ();
 sky130_fd_sc_hd__nand2_1 _17994_ (.A(\cs_registers_i.dscratch0_q[17] ),
    .B(_12315_),
    .Y(_12327_));
 sky130_fd_sc_hd__o21ai_0 _17995_ (.A1(_11294_),
    .A2(_12315_),
    .B1(_12327_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _17996_ (.A(\cs_registers_i.dscratch0_q[18] ),
    .B(_12315_),
    .Y(_12328_));
 sky130_fd_sc_hd__o21ai_0 _17997_ (.A1(_11319_),
    .A2(_12315_),
    .B1(_12328_),
    .Y(_00197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_728 ();
 sky130_fd_sc_hd__nand2_1 _17999_ (.A(\cs_registers_i.dscratch0_q[19] ),
    .B(_12315_),
    .Y(_12330_));
 sky130_fd_sc_hd__o21ai_0 _18000_ (.A1(_11333_),
    .A2(_12315_),
    .B1(_12330_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _18001_ (.A(\cs_registers_i.dscratch0_q[1] ),
    .B(_12315_),
    .Y(_12331_));
 sky130_fd_sc_hd__o21ai_0 _18002_ (.A1(_11354_),
    .A2(_12315_),
    .B1(_12331_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _18003_ (.A(\cs_registers_i.dscratch0_q[20] ),
    .B(_12315_),
    .Y(_12332_));
 sky130_fd_sc_hd__o21ai_0 _18004_ (.A1(_11369_),
    .A2(_12315_),
    .B1(_12332_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _18005_ (.A(\cs_registers_i.dscratch0_q[21] ),
    .B(_12315_),
    .Y(_12333_));
 sky130_fd_sc_hd__o21ai_0 _18006_ (.A1(_11390_),
    .A2(_12315_),
    .B1(_12333_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _18007_ (.A(\cs_registers_i.dscratch0_q[22] ),
    .B(_12315_),
    .Y(_12334_));
 sky130_fd_sc_hd__o21ai_0 _18008_ (.A1(_11406_),
    .A2(_12315_),
    .B1(_12334_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _18009_ (.A(\cs_registers_i.dscratch0_q[23] ),
    .B(_12315_),
    .Y(_12335_));
 sky130_fd_sc_hd__o21ai_0 _18010_ (.A1(_11426_),
    .A2(_12315_),
    .B1(_12335_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _18011_ (.A(\cs_registers_i.dscratch0_q[24] ),
    .B(_12315_),
    .Y(_12336_));
 sky130_fd_sc_hd__o21ai_0 _18012_ (.A1(_11441_),
    .A2(_12315_),
    .B1(_12336_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _18013_ (.A(\cs_registers_i.dscratch0_q[25] ),
    .B(_12315_),
    .Y(_12337_));
 sky130_fd_sc_hd__o21ai_0 _18014_ (.A1(_11457_),
    .A2(_12315_),
    .B1(_12337_),
    .Y(_00205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_727 ();
 sky130_fd_sc_hd__nand2_1 _18016_ (.A(\cs_registers_i.dscratch0_q[26] ),
    .B(_12315_),
    .Y(_12339_));
 sky130_fd_sc_hd__o21ai_0 _18017_ (.A1(_11476_),
    .A2(_12315_),
    .B1(_12339_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _18018_ (.A(\cs_registers_i.dscratch0_q[27] ),
    .B(_12315_),
    .Y(_12340_));
 sky130_fd_sc_hd__o21ai_0 _18019_ (.A1(_11490_),
    .A2(_12315_),
    .B1(_12340_),
    .Y(_00207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_726 ();
 sky130_fd_sc_hd__nand2_1 _18021_ (.A(\cs_registers_i.dscratch0_q[28] ),
    .B(_12315_),
    .Y(_12342_));
 sky130_fd_sc_hd__o21ai_0 _18022_ (.A1(net3480),
    .A2(_12315_),
    .B1(_12342_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _18023_ (.A(\cs_registers_i.dscratch0_q[29] ),
    .B(_12315_),
    .Y(_12343_));
 sky130_fd_sc_hd__o21ai_0 _18024_ (.A1(_11530_),
    .A2(_12315_),
    .B1(_12343_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _18025_ (.A(\cs_registers_i.dscratch0_q[2] ),
    .B(_12315_),
    .Y(_12344_));
 sky130_fd_sc_hd__o21ai_0 _18026_ (.A1(_11082_),
    .A2(_12315_),
    .B1(_12344_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _18027_ (.A(\cs_registers_i.dscratch0_q[30] ),
    .B(_12315_),
    .Y(_12345_));
 sky130_fd_sc_hd__o21ai_0 _18028_ (.A1(_11550_),
    .A2(_12315_),
    .B1(_12345_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _18029_ (.A(\cs_registers_i.dscratch0_q[31] ),
    .B(_12315_),
    .Y(_12346_));
 sky130_fd_sc_hd__o21ai_0 _18030_ (.A1(_11565_),
    .A2(_12315_),
    .B1(_12346_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(\cs_registers_i.dscratch0_q[3] ),
    .B(_12315_),
    .Y(_12347_));
 sky130_fd_sc_hd__o21ai_0 _18032_ (.A1(_11612_),
    .A2(_12315_),
    .B1(_12347_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _18033_ (.A(\cs_registers_i.dscratch0_q[4] ),
    .B(_12315_),
    .Y(_12348_));
 sky130_fd_sc_hd__o21ai_0 _18034_ (.A1(_11780_),
    .A2(_12315_),
    .B1(_12348_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _18035_ (.A(\cs_registers_i.dscratch0_q[5] ),
    .B(_12315_),
    .Y(_12349_));
 sky130_fd_sc_hd__o21ai_0 _18036_ (.A1(_11647_),
    .A2(_12315_),
    .B1(_12349_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _18037_ (.A(\cs_registers_i.dscratch0_q[6] ),
    .B(_12315_),
    .Y(_12350_));
 sky130_fd_sc_hd__o21ai_0 _18038_ (.A1(_11664_),
    .A2(_12315_),
    .B1(_12350_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _18039_ (.A(\cs_registers_i.dscratch0_q[7] ),
    .B(_12315_),
    .Y(_12351_));
 sky130_fd_sc_hd__o21ai_0 _18040_ (.A1(net3478),
    .A2(_12315_),
    .B1(_12351_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _18041_ (.A(\cs_registers_i.dscratch0_q[8] ),
    .B(_12315_),
    .Y(_12352_));
 sky130_fd_sc_hd__o21ai_0 _18042_ (.A1(_11707_),
    .A2(_12315_),
    .B1(_12352_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(\cs_registers_i.dscratch0_q[9] ),
    .B(_12315_),
    .Y(_12353_));
 sky130_fd_sc_hd__o21ai_0 _18044_ (.A1(_11726_),
    .A2(_12315_),
    .B1(_12353_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_8 _18045_ (.A(net3501),
    .B(_11227_),
    .Y(_12354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_724 ();
 sky130_fd_sc_hd__nand2_1 _18048_ (.A(\cs_registers_i.dscratch1_q[0] ),
    .B(_12354_),
    .Y(_12357_));
 sky130_fd_sc_hd__o21ai_0 _18049_ (.A1(_11042_),
    .A2(_12354_),
    .B1(_12357_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _18050_ (.A(\cs_registers_i.dscratch1_q[10] ),
    .B(_12354_),
    .Y(_12358_));
 sky130_fd_sc_hd__o21ai_0 _18051_ (.A1(_11145_),
    .A2(_12354_),
    .B1(_12358_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _18052_ (.A(\cs_registers_i.dscratch1_q[11] ),
    .B(_12354_),
    .Y(_12359_));
 sky130_fd_sc_hd__o21ai_0 _18053_ (.A1(_11177_),
    .A2(_12354_),
    .B1(_12359_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _18054_ (.A(\cs_registers_i.dscratch1_q[12] ),
    .B(_12354_),
    .Y(_12360_));
 sky130_fd_sc_hd__o21ai_0 _18055_ (.A1(_11197_),
    .A2(_12354_),
    .B1(_12360_),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(\cs_registers_i.dscratch1_q[13] ),
    .B(_12354_),
    .Y(_12361_));
 sky130_fd_sc_hd__o21ai_0 _18057_ (.A1(_11214_),
    .A2(_12354_),
    .B1(_12361_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _18058_ (.A(\cs_registers_i.dscratch1_q[14] ),
    .B(_12354_),
    .Y(_12362_));
 sky130_fd_sc_hd__o21ai_0 _18059_ (.A1(_11235_),
    .A2(_12354_),
    .B1(_12362_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _18060_ (.A(\cs_registers_i.dscratch1_q[15] ),
    .B(_12354_),
    .Y(_12363_));
 sky130_fd_sc_hd__o21ai_0 _18061_ (.A1(_11255_),
    .A2(_12354_),
    .B1(_12363_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _18062_ (.A(\cs_registers_i.dscratch1_q[16] ),
    .B(_12354_),
    .Y(_12364_));
 sky130_fd_sc_hd__o21ai_0 _18063_ (.A1(_11270_),
    .A2(_12354_),
    .B1(_12364_),
    .Y(_00227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_723 ();
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(\cs_registers_i.dscratch1_q[17] ),
    .B(_12354_),
    .Y(_12366_));
 sky130_fd_sc_hd__o21ai_0 _18066_ (.A1(_11294_),
    .A2(_12354_),
    .B1(_12366_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _18067_ (.A(\cs_registers_i.dscratch1_q[18] ),
    .B(_12354_),
    .Y(_12367_));
 sky130_fd_sc_hd__o21ai_0 _18068_ (.A1(_11319_),
    .A2(_12354_),
    .B1(_12367_),
    .Y(_00229_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_722 ();
 sky130_fd_sc_hd__nand2_1 _18070_ (.A(\cs_registers_i.dscratch1_q[19] ),
    .B(_12354_),
    .Y(_12369_));
 sky130_fd_sc_hd__o21ai_0 _18071_ (.A1(_11333_),
    .A2(_12354_),
    .B1(_12369_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(\cs_registers_i.dscratch1_q[1] ),
    .B(_12354_),
    .Y(_12370_));
 sky130_fd_sc_hd__o21ai_0 _18073_ (.A1(_11354_),
    .A2(_12354_),
    .B1(_12370_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _18074_ (.A(\cs_registers_i.dscratch1_q[20] ),
    .B(_12354_),
    .Y(_12371_));
 sky130_fd_sc_hd__o21ai_0 _18075_ (.A1(_11369_),
    .A2(_12354_),
    .B1(_12371_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _18076_ (.A(\cs_registers_i.dscratch1_q[21] ),
    .B(_12354_),
    .Y(_12372_));
 sky130_fd_sc_hd__o21ai_0 _18077_ (.A1(_11390_),
    .A2(_12354_),
    .B1(_12372_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _18078_ (.A(\cs_registers_i.dscratch1_q[22] ),
    .B(_12354_),
    .Y(_12373_));
 sky130_fd_sc_hd__o21ai_0 _18079_ (.A1(_11406_),
    .A2(_12354_),
    .B1(_12373_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _18080_ (.A(\cs_registers_i.dscratch1_q[23] ),
    .B(_12354_),
    .Y(_12374_));
 sky130_fd_sc_hd__o21ai_0 _18081_ (.A1(net3492),
    .A2(_12354_),
    .B1(_12374_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(\cs_registers_i.dscratch1_q[24] ),
    .B(_12354_),
    .Y(_12375_));
 sky130_fd_sc_hd__o21ai_0 _18083_ (.A1(_11441_),
    .A2(_12354_),
    .B1(_12375_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _18084_ (.A(\cs_registers_i.dscratch1_q[25] ),
    .B(_12354_),
    .Y(_12376_));
 sky130_fd_sc_hd__o21ai_0 _18085_ (.A1(_11457_),
    .A2(_12354_),
    .B1(_12376_),
    .Y(_00237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_721 ();
 sky130_fd_sc_hd__nand2_1 _18087_ (.A(\cs_registers_i.dscratch1_q[26] ),
    .B(_12354_),
    .Y(_12378_));
 sky130_fd_sc_hd__o21ai_0 _18088_ (.A1(_11476_),
    .A2(_12354_),
    .B1(_12378_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _18089_ (.A(\cs_registers_i.dscratch1_q[27] ),
    .B(_12354_),
    .Y(_12379_));
 sky130_fd_sc_hd__o21ai_0 _18090_ (.A1(_11490_),
    .A2(_12354_),
    .B1(_12379_),
    .Y(_00239_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_720 ();
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(\cs_registers_i.dscratch1_q[28] ),
    .B(_12354_),
    .Y(_12381_));
 sky130_fd_sc_hd__o21ai_0 _18093_ (.A1(net3480),
    .A2(_12354_),
    .B1(_12381_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _18094_ (.A(\cs_registers_i.dscratch1_q[29] ),
    .B(_12354_),
    .Y(_12382_));
 sky130_fd_sc_hd__o21ai_0 _18095_ (.A1(_11530_),
    .A2(_12354_),
    .B1(_12382_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _18096_ (.A(\cs_registers_i.dscratch1_q[2] ),
    .B(_12354_),
    .Y(_12383_));
 sky130_fd_sc_hd__o21ai_0 _18097_ (.A1(_11082_),
    .A2(_12354_),
    .B1(_12383_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _18098_ (.A(\cs_registers_i.dscratch1_q[30] ),
    .B(_12354_),
    .Y(_12384_));
 sky130_fd_sc_hd__o21ai_0 _18099_ (.A1(_11550_),
    .A2(_12354_),
    .B1(_12384_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _18100_ (.A(\cs_registers_i.dscratch1_q[31] ),
    .B(_12354_),
    .Y(_12385_));
 sky130_fd_sc_hd__o21ai_0 _18101_ (.A1(_11565_),
    .A2(_12354_),
    .B1(_12385_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(\cs_registers_i.dscratch1_q[3] ),
    .B(_12354_),
    .Y(_12386_));
 sky130_fd_sc_hd__o21ai_0 _18103_ (.A1(_11612_),
    .A2(_12354_),
    .B1(_12386_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(\cs_registers_i.dscratch1_q[4] ),
    .B(_12354_),
    .Y(_12387_));
 sky130_fd_sc_hd__o21ai_0 _18105_ (.A1(_11780_),
    .A2(_12354_),
    .B1(_12387_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _18106_ (.A(\cs_registers_i.dscratch1_q[5] ),
    .B(_12354_),
    .Y(_12388_));
 sky130_fd_sc_hd__o21ai_0 _18107_ (.A1(_11647_),
    .A2(_12354_),
    .B1(_12388_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _18108_ (.A(\cs_registers_i.dscratch1_q[6] ),
    .B(_12354_),
    .Y(_12389_));
 sky130_fd_sc_hd__o21ai_0 _18109_ (.A1(_11664_),
    .A2(_12354_),
    .B1(_12389_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _18110_ (.A(\cs_registers_i.dscratch1_q[7] ),
    .B(_12354_),
    .Y(_12390_));
 sky130_fd_sc_hd__o21ai_0 _18111_ (.A1(_11685_),
    .A2(_12354_),
    .B1(_12390_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _18112_ (.A(\cs_registers_i.dscratch1_q[8] ),
    .B(_12354_),
    .Y(_12391_));
 sky130_fd_sc_hd__o21ai_0 _18113_ (.A1(_11707_),
    .A2(_12354_),
    .B1(_12391_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _18114_ (.A(\cs_registers_i.dscratch1_q[9] ),
    .B(_12354_),
    .Y(_12392_));
 sky130_fd_sc_hd__o21ai_0 _18115_ (.A1(_11726_),
    .A2(_12354_),
    .B1(_12392_),
    .Y(_00251_));
 sky130_fd_sc_hd__nor2_4 _18116_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_12188_),
    .Y(_12393_));
 sky130_fd_sc_hd__and2_4 _18117_ (.A(net3545),
    .B(_12393_),
    .X(_12394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_719 ();
 sky130_fd_sc_hd__nor4_4 _18119_ (.A(_10500_),
    .B(_10505_),
    .C(_10512_),
    .D(_10784_),
    .Y(_12396_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_716 ();
 sky130_fd_sc_hd__and2_4 _18123_ (.A(\cs_registers_i.nmi_mode_i ),
    .B(net3663),
    .X(_12400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_715 ();
 sky130_fd_sc_hd__nor2_4 _18125_ (.A(_12394_),
    .B(_12400_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_4 _18126_ (.A(_10613_),
    .B(net3501),
    .Y(_12403_));
 sky130_fd_sc_hd__nand2_8 _18127_ (.A(_12402_),
    .B(_12403_),
    .Y(_12404_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_714 ();
 sky130_fd_sc_hd__or2_4 _18129_ (.A(_12394_),
    .B(_12400_),
    .X(_12406_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_713 ();
 sky130_fd_sc_hd__nor2_2 _18131_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.load_err_q ),
    .Y(_12408_));
 sky130_fd_sc_hd__nor2_1 _18132_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10648_),
    .Y(_12409_));
 sky130_fd_sc_hd__a21oi_2 _18133_ (.A1(_12408_),
    .A2(_12409_),
    .B1(_12168_),
    .Y(_12410_));
 sky130_fd_sc_hd__nor2_1 _18134_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10647_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand3_1 _18135_ (.A(net3895),
    .B(_10646_),
    .C(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__or3_4 _18136_ (.A(net3895),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .C(_10787_),
    .X(_12413_));
 sky130_fd_sc_hd__nand2_1 _18137_ (.A(\cs_registers_i.priv_mode_id_o[1] ),
    .B(net3950),
    .Y(_12414_));
 sky130_fd_sc_hd__o32a_1 _18138_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10791_),
    .A3(_12412_),
    .B1(_12413_),
    .B2(_12414_),
    .X(_12415_));
 sky130_fd_sc_hd__and2_4 _18139_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .X(_12416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_712 ();
 sky130_fd_sc_hd__nor3_2 _18141_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10648_),
    .C(_12408_),
    .Y(_12418_));
 sky130_fd_sc_hd__nor2_1 _18142_ (.A(_12416_),
    .B(_12418_),
    .Y(_12419_));
 sky130_fd_sc_hd__nand2_2 _18143_ (.A(_12415_),
    .B(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(\cs_registers_i.mie_q[10] ),
    .B(net131),
    .Y(_12421_));
 sky130_fd_sc_hd__nand2_1 _18145_ (.A(\cs_registers_i.mie_q[2] ),
    .B(net137),
    .Y(_12422_));
 sky130_fd_sc_hd__a32oi_1 _18146_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net136),
    .A3(_12422_),
    .B1(net138),
    .B2(\cs_registers_i.mie_q[3] ),
    .Y(_12423_));
 sky130_fd_sc_hd__a21oi_1 _18147_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net139),
    .B1(_12423_),
    .Y(_12424_));
 sky130_fd_sc_hd__a21oi_2 _18148_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net140),
    .B1(_12424_),
    .Y(_12425_));
 sky130_fd_sc_hd__a21oi_1 _18149_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net141),
    .B1(_12425_),
    .Y(_12426_));
 sky130_fd_sc_hd__a21oi_2 _18150_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net142),
    .B1(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__nand2_1 _18151_ (.A(\cs_registers_i.mie_q[9] ),
    .B(net144),
    .Y(_12428_));
 sky130_fd_sc_hd__o21ai_4 _18152_ (.A1(_10813_),
    .A2(_12427_),
    .B1(_12428_),
    .Y(_12429_));
 sky130_fd_sc_hd__a22o_1 _18153_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(net132),
    .B1(_12421_),
    .B2(_12429_),
    .X(_12430_));
 sky130_fd_sc_hd__a22o_1 _18154_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(net134),
    .B1(_10810_),
    .B2(_12430_),
    .X(_12431_));
 sky130_fd_sc_hd__a221oi_2 _18155_ (.A1(_10822_),
    .A2(net145),
    .B1(_10816_),
    .B2(_12431_),
    .C1(_10817_),
    .Y(_12432_));
 sky130_fd_sc_hd__nor2b_4 _18156_ (.A(_12432_),
    .B_N(_12170_),
    .Y(_12433_));
 sky130_fd_sc_hd__a21oi_4 _18157_ (.A1(_12410_),
    .A2(_12420_),
    .B1(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__nand2_8 _18158_ (.A(net3545),
    .B(_12393_),
    .Y(_12435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_710 ();
 sky130_fd_sc_hd__nand2_1 _18161_ (.A(\cs_registers_i.mstack_cause_q[0] ),
    .B(_12400_),
    .Y(_12438_));
 sky130_fd_sc_hd__o221a_1 _18162_ (.A1(_11042_),
    .A2(_12406_),
    .B1(_12434_),
    .B2(_12435_),
    .C1(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__nor2_1 _18163_ (.A(\cs_registers_i.mcause_q[0] ),
    .B(_12404_),
    .Y(_12440_));
 sky130_fd_sc_hd__a21oi_1 _18164_ (.A1(_12404_),
    .A2(_12439_),
    .B1(_12440_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2b_1 _18165_ (.A_N(_11354_),
    .B(_12402_),
    .Y(_12441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_708 ();
 sky130_fd_sc_hd__o21ai_2 _18168_ (.A1(_10804_),
    .A2(_10807_),
    .B1(_10805_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand2_4 _18169_ (.A(_10814_),
    .B(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_2 _18170_ (.A(_10810_),
    .B(_10811_),
    .Y(_12446_));
 sky130_fd_sc_hd__a21oi_2 _18171_ (.A1(_10812_),
    .A2(_12445_),
    .B1(_12446_),
    .Y(_12447_));
 sky130_fd_sc_hd__nand2_4 _18172_ (.A(_10822_),
    .B(net145),
    .Y(_12448_));
 sky130_fd_sc_hd__nand2_4 _18173_ (.A(_10816_),
    .B(_12448_),
    .Y(_12449_));
 sky130_fd_sc_hd__o31ai_4 _18174_ (.A1(_10817_),
    .A2(_12447_),
    .A3(_12449_),
    .B1(_12170_),
    .Y(_12450_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_707 ();
 sky130_fd_sc_hd__and2_4 _18176_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10646_),
    .X(_12452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_706 ();
 sky130_fd_sc_hd__a31oi_1 _18178_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(_10646_),
    .A3(_10647_),
    .B1(_12452_),
    .Y(_12454_));
 sky130_fd_sc_hd__nand2_1 _18179_ (.A(_12415_),
    .B(_12454_),
    .Y(_12455_));
 sky130_fd_sc_hd__nand2_1 _18180_ (.A(_12410_),
    .B(_12455_),
    .Y(_12456_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_705 ();
 sky130_fd_sc_hd__a21oi_1 _18182_ (.A1(_12450_),
    .A2(_12456_),
    .B1(_12435_),
    .Y(_12458_));
 sky130_fd_sc_hd__a21oi_1 _18183_ (.A1(\cs_registers_i.mstack_cause_q[1] ),
    .A2(_12400_),
    .B1(_12458_),
    .Y(_12459_));
 sky130_fd_sc_hd__nor2_1 _18184_ (.A(\cs_registers_i.mcause_q[1] ),
    .B(_12404_),
    .Y(_12460_));
 sky130_fd_sc_hd__a31oi_1 _18185_ (.A1(_12404_),
    .A2(_12441_),
    .A3(_12459_),
    .B1(_12460_),
    .Y(_00253_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_704 ();
 sky130_fd_sc_hd__nor2_1 _18187_ (.A(_11082_),
    .B(_12406_),
    .Y(_12462_));
 sky130_fd_sc_hd__nand2_1 _18188_ (.A(_10812_),
    .B(_10814_),
    .Y(_12463_));
 sky130_fd_sc_hd__nor2_2 _18189_ (.A(_10806_),
    .B(_12463_),
    .Y(_12464_));
 sky130_fd_sc_hd__o41ai_4 _18190_ (.A1(_12446_),
    .A2(_10820_),
    .A3(_12449_),
    .A4(_12464_),
    .B1(_12170_),
    .Y(_12465_));
 sky130_fd_sc_hd__nand2_1 _18191_ (.A(_10783_),
    .B(_12418_),
    .Y(_12466_));
 sky130_fd_sc_hd__a21oi_1 _18192_ (.A1(_12465_),
    .A2(_12466_),
    .B1(_12435_),
    .Y(_12467_));
 sky130_fd_sc_hd__a211oi_1 _18193_ (.A1(\cs_registers_i.mstack_cause_q[2] ),
    .A2(_12400_),
    .B1(_12462_),
    .C1(_12467_),
    .Y(_12468_));
 sky130_fd_sc_hd__nor2_1 _18194_ (.A(\cs_registers_i.mcause_q[2] ),
    .B(_12404_),
    .Y(_12469_));
 sky130_fd_sc_hd__a21oi_1 _18195_ (.A1(_12404_),
    .A2(_12468_),
    .B1(_12469_),
    .Y(_00254_));
 sky130_fd_sc_hd__nor2_1 _18196_ (.A(_10809_),
    .B(_10818_),
    .Y(_12470_));
 sky130_fd_sc_hd__o31ai_4 _18197_ (.A1(_10815_),
    .A2(_12449_),
    .A3(_12470_),
    .B1(_12170_),
    .Y(_12471_));
 sky130_fd_sc_hd__o21ai_2 _18198_ (.A1(_12168_),
    .A2(_12413_),
    .B1(_12471_),
    .Y(_12472_));
 sky130_fd_sc_hd__nand2_1 _18199_ (.A(_12393_),
    .B(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__o21ai_0 _18200_ (.A1(_11612_),
    .A2(_12393_),
    .B1(_12473_),
    .Y(_12474_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_703 ();
 sky130_fd_sc_hd__nor2_1 _18202_ (.A(net3545),
    .B(net3663),
    .Y(_12476_));
 sky130_fd_sc_hd__a21oi_1 _18203_ (.A1(_10822_),
    .A2(net3663),
    .B1(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__nor2_1 _18204_ (.A(_11612_),
    .B(_12477_),
    .Y(_12478_));
 sky130_fd_sc_hd__a221oi_1 _18205_ (.A1(\cs_registers_i.mstack_cause_q[3] ),
    .A2(_12400_),
    .B1(_12474_),
    .B2(net3545),
    .C1(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__nor2_1 _18206_ (.A(\cs_registers_i.mcause_q[3] ),
    .B(_12404_),
    .Y(_12480_));
 sky130_fd_sc_hd__a21oi_1 _18207_ (.A1(_12404_),
    .A2(_12479_),
    .B1(_12480_),
    .Y(_00255_));
 sky130_fd_sc_hd__a21boi_4 _18208_ (.A1(_10817_),
    .A2(_12448_),
    .B1_N(net3573),
    .Y(_12481_));
 sky130_fd_sc_hd__a221oi_1 _18209_ (.A1(\cs_registers_i.mstack_cause_q[4] ),
    .A2(_12400_),
    .B1(_12402_),
    .B2(_11631_),
    .C1(_12481_),
    .Y(_12482_));
 sky130_fd_sc_hd__nor2_1 _18210_ (.A(\cs_registers_i.mcause_q[4] ),
    .B(_12404_),
    .Y(_12483_));
 sky130_fd_sc_hd__a21oi_1 _18211_ (.A1(_12404_),
    .A2(_12482_),
    .B1(_12483_),
    .Y(_00256_));
 sky130_fd_sc_hd__nor2_1 _18212_ (.A(_11565_),
    .B(_12406_),
    .Y(_12484_));
 sky130_fd_sc_hd__a211oi_1 _18213_ (.A1(\cs_registers_i.mstack_cause_q[5] ),
    .A2(_12400_),
    .B1(_12484_),
    .C1(net3573),
    .Y(_12485_));
 sky130_fd_sc_hd__nor2_1 _18214_ (.A(\cs_registers_i.mcause_q[5] ),
    .B(_12404_),
    .Y(_12486_));
 sky130_fd_sc_hd__a21oi_1 _18215_ (.A1(_12404_),
    .A2(_12485_),
    .B1(_12486_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_4 _18216_ (.A(net3538),
    .B(net3501),
    .Y(_12487_));
 sky130_fd_sc_hd__a32o_1 _18217_ (.A1(\cs_registers_i.csr_mepc_o[0] ),
    .A2(_12402_),
    .A3(_12487_),
    .B1(\cs_registers_i.mstack_epc_q[0] ),
    .B2(_12400_),
    .X(_00258_));
 sky130_fd_sc_hd__nand2_8 _18218_ (.A(_12402_),
    .B(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_702 ();
 sky130_fd_sc_hd__nand2_1 _18220_ (.A(\cs_registers_i.mstack_epc_q[10] ),
    .B(_12400_),
    .Y(_12490_));
 sky130_fd_sc_hd__o221a_1 _18221_ (.A1(_12207_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11145_),
    .C1(_12490_),
    .X(_12491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_701 ();
 sky130_fd_sc_hd__nor2_1 _18223_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(_12488_),
    .Y(_12493_));
 sky130_fd_sc_hd__a21oi_1 _18224_ (.A1(_12488_),
    .A2(_12491_),
    .B1(_12493_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _18225_ (.A(\cs_registers_i.mstack_epc_q[11] ),
    .B(_12400_),
    .Y(_12494_));
 sky130_fd_sc_hd__o221a_1 _18226_ (.A1(_12213_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11177_),
    .C1(_12494_),
    .X(_12495_));
 sky130_fd_sc_hd__nor2_1 _18227_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(_12488_),
    .Y(_12496_));
 sky130_fd_sc_hd__a21oi_1 _18228_ (.A1(_12488_),
    .A2(_12495_),
    .B1(_12496_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _18229_ (.A(\cs_registers_i.mstack_epc_q[12] ),
    .B(_12400_),
    .Y(_12497_));
 sky130_fd_sc_hd__o221a_1 _18230_ (.A1(_12216_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11197_),
    .C1(_12497_),
    .X(_12498_));
 sky130_fd_sc_hd__nor2_1 _18231_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(_12488_),
    .Y(_12499_));
 sky130_fd_sc_hd__a21oi_1 _18232_ (.A1(_12488_),
    .A2(_12498_),
    .B1(_12499_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _18233_ (.A(\cs_registers_i.mstack_epc_q[13] ),
    .B(_12400_),
    .Y(_12500_));
 sky130_fd_sc_hd__o221a_1 _18234_ (.A1(_12219_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11214_),
    .C1(_12500_),
    .X(_12501_));
 sky130_fd_sc_hd__nor2_1 _18235_ (.A(\cs_registers_i.csr_mepc_o[13] ),
    .B(_12488_),
    .Y(_12502_));
 sky130_fd_sc_hd__a21oi_1 _18236_ (.A1(_12488_),
    .A2(_12501_),
    .B1(_12502_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _18237_ (.A(\cs_registers_i.mstack_epc_q[14] ),
    .B(_12400_),
    .Y(_12503_));
 sky130_fd_sc_hd__o221a_1 _18238_ (.A1(_12222_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11235_),
    .C1(_12503_),
    .X(_12504_));
 sky130_fd_sc_hd__nor2_1 _18239_ (.A(\cs_registers_i.csr_mepc_o[14] ),
    .B(_12488_),
    .Y(_12505_));
 sky130_fd_sc_hd__a21oi_1 _18240_ (.A1(_12488_),
    .A2(_12504_),
    .B1(_12505_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _18241_ (.A(\cs_registers_i.mstack_epc_q[15] ),
    .B(_12400_),
    .Y(_12506_));
 sky130_fd_sc_hd__o221a_1 _18242_ (.A1(_12227_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11255_),
    .C1(_12506_),
    .X(_12507_));
 sky130_fd_sc_hd__nor2_1 _18243_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(_12488_),
    .Y(_12508_));
 sky130_fd_sc_hd__a21oi_1 _18244_ (.A1(_12488_),
    .A2(_12507_),
    .B1(_12508_),
    .Y(_00264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_700 ();
 sky130_fd_sc_hd__nand2_1 _18246_ (.A(\cs_registers_i.mstack_epc_q[16] ),
    .B(_12400_),
    .Y(_12510_));
 sky130_fd_sc_hd__o221a_1 _18247_ (.A1(_12230_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11270_),
    .C1(_12510_),
    .X(_12511_));
 sky130_fd_sc_hd__nor2_1 _18248_ (.A(\cs_registers_i.csr_mepc_o[16] ),
    .B(_12488_),
    .Y(_12512_));
 sky130_fd_sc_hd__a21oi_1 _18249_ (.A1(_12488_),
    .A2(_12511_),
    .B1(_12512_),
    .Y(_00265_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_698 ();
 sky130_fd_sc_hd__nand2_1 _18252_ (.A(\cs_registers_i.mstack_epc_q[17] ),
    .B(_12400_),
    .Y(_12515_));
 sky130_fd_sc_hd__o221a_1 _18253_ (.A1(_12233_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11294_),
    .C1(_12515_),
    .X(_12516_));
 sky130_fd_sc_hd__nor2_1 _18254_ (.A(\cs_registers_i.csr_mepc_o[17] ),
    .B(_12488_),
    .Y(_12517_));
 sky130_fd_sc_hd__a21oi_1 _18255_ (.A1(_12488_),
    .A2(_12516_),
    .B1(_12517_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _18256_ (.A(\cs_registers_i.mstack_epc_q[18] ),
    .B(_12400_),
    .Y(_12518_));
 sky130_fd_sc_hd__o221a_1 _18257_ (.A1(_12236_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11319_),
    .C1(_12518_),
    .X(_12519_));
 sky130_fd_sc_hd__nor2_1 _18258_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(_12488_),
    .Y(_12520_));
 sky130_fd_sc_hd__a21oi_1 _18259_ (.A1(_12488_),
    .A2(_12519_),
    .B1(_12520_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _18260_ (.A(\cs_registers_i.mstack_epc_q[19] ),
    .B(_12400_),
    .Y(_12521_));
 sky130_fd_sc_hd__o221a_1 _18261_ (.A1(_12239_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11333_),
    .C1(_12521_),
    .X(_12522_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_697 ();
 sky130_fd_sc_hd__nor2_1 _18263_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(_12488_),
    .Y(_12524_));
 sky130_fd_sc_hd__a21oi_1 _18264_ (.A1(_12488_),
    .A2(_12522_),
    .B1(_12524_),
    .Y(_00268_));
 sky130_fd_sc_hd__nor2_1 _18265_ (.A(_12246_),
    .B(_12435_),
    .Y(_12525_));
 sky130_fd_sc_hd__a21oi_1 _18266_ (.A1(\cs_registers_i.mstack_epc_q[1] ),
    .A2(_12400_),
    .B1(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nor2_1 _18267_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(_12488_),
    .Y(_12527_));
 sky130_fd_sc_hd__a31oi_1 _18268_ (.A1(_12441_),
    .A2(_12488_),
    .A3(_12526_),
    .B1(_12527_),
    .Y(_00269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_696 ();
 sky130_fd_sc_hd__nand2_1 _18270_ (.A(\cs_registers_i.mstack_epc_q[20] ),
    .B(_12400_),
    .Y(_12529_));
 sky130_fd_sc_hd__o221a_1 _18271_ (.A1(_12250_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11369_),
    .C1(_12529_),
    .X(_12530_));
 sky130_fd_sc_hd__nor2_1 _18272_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(_12488_),
    .Y(_12531_));
 sky130_fd_sc_hd__a21oi_1 _18273_ (.A1(_12488_),
    .A2(_12530_),
    .B1(_12531_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _18274_ (.A(\cs_registers_i.mstack_epc_q[21] ),
    .B(_12400_),
    .Y(_12532_));
 sky130_fd_sc_hd__o221a_1 _18275_ (.A1(_12253_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11390_),
    .C1(_12532_),
    .X(_12533_));
 sky130_fd_sc_hd__nor2_1 _18276_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(_12488_),
    .Y(_12534_));
 sky130_fd_sc_hd__a21oi_1 _18277_ (.A1(_12488_),
    .A2(_12533_),
    .B1(_12534_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _18278_ (.A(\cs_registers_i.mstack_epc_q[22] ),
    .B(_12400_),
    .Y(_12535_));
 sky130_fd_sc_hd__o221a_1 _18279_ (.A1(_12256_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11406_),
    .C1(_12535_),
    .X(_12536_));
 sky130_fd_sc_hd__nor2_1 _18280_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(_12488_),
    .Y(_12537_));
 sky130_fd_sc_hd__a21oi_1 _18281_ (.A1(_12488_),
    .A2(_12536_),
    .B1(_12537_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _18282_ (.A(\cs_registers_i.mstack_epc_q[23] ),
    .B(_12400_),
    .Y(_12538_));
 sky130_fd_sc_hd__o221a_1 _18283_ (.A1(_12259_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11426_),
    .C1(_12538_),
    .X(_12539_));
 sky130_fd_sc_hd__nor2_1 _18284_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(_12488_),
    .Y(_12540_));
 sky130_fd_sc_hd__a21oi_1 _18285_ (.A1(_12488_),
    .A2(_12539_),
    .B1(_12540_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _18286_ (.A(_10822_),
    .B(_11441_),
    .Y(_12541_));
 sky130_fd_sc_hd__o22ai_1 _18287_ (.A1(_12263_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11441_),
    .Y(_12542_));
 sky130_fd_sc_hd__a31oi_1 _18288_ (.A1(\cs_registers_i.mstack_epc_q[24] ),
    .A2(net3663),
    .A3(_12541_),
    .B1(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(_12488_),
    .Y(_12544_));
 sky130_fd_sc_hd__a21oi_1 _18290_ (.A1(_12488_),
    .A2(_12543_),
    .B1(_12544_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _18291_ (.A(\cs_registers_i.mstack_epc_q[25] ),
    .B(_12400_),
    .Y(_12545_));
 sky130_fd_sc_hd__o221a_1 _18292_ (.A1(_12266_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11457_),
    .C1(_12545_),
    .X(_12546_));
 sky130_fd_sc_hd__nor2_1 _18293_ (.A(\cs_registers_i.csr_mepc_o[25] ),
    .B(_12488_),
    .Y(_12547_));
 sky130_fd_sc_hd__a21oi_1 _18294_ (.A1(_12488_),
    .A2(_12546_),
    .B1(_12547_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _18295_ (.A(\cs_registers_i.mstack_epc_q[26] ),
    .B(_12400_),
    .Y(_12548_));
 sky130_fd_sc_hd__o221a_1 _18296_ (.A1(_12270_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11476_),
    .C1(_12548_),
    .X(_12549_));
 sky130_fd_sc_hd__nor2_1 _18297_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(_12488_),
    .Y(_12550_));
 sky130_fd_sc_hd__a21oi_1 _18298_ (.A1(_12488_),
    .A2(_12549_),
    .B1(_12550_),
    .Y(_00276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_695 ();
 sky130_fd_sc_hd__nand2_1 _18300_ (.A(\cs_registers_i.mstack_epc_q[27] ),
    .B(_12400_),
    .Y(_12552_));
 sky130_fd_sc_hd__o221a_1 _18301_ (.A1(_12273_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11490_),
    .C1(_12552_),
    .X(_12553_));
 sky130_fd_sc_hd__nor2_1 _18302_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(_12488_),
    .Y(_12554_));
 sky130_fd_sc_hd__a21oi_1 _18303_ (.A1(_12488_),
    .A2(_12553_),
    .B1(_12554_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(\cs_registers_i.mstack_epc_q[28] ),
    .B(_12400_),
    .Y(_12555_));
 sky130_fd_sc_hd__o221a_1 _18305_ (.A1(_12276_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11506_),
    .C1(_12555_),
    .X(_12556_));
 sky130_fd_sc_hd__nor2_1 _18306_ (.A(\cs_registers_i.csr_mepc_o[28] ),
    .B(_12488_),
    .Y(_12557_));
 sky130_fd_sc_hd__a21oi_1 _18307_ (.A1(_12488_),
    .A2(_12556_),
    .B1(_12557_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _18308_ (.A(\cs_registers_i.mstack_epc_q[29] ),
    .B(_12400_),
    .Y(_12558_));
 sky130_fd_sc_hd__o221a_1 _18309_ (.A1(_12281_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11530_),
    .C1(_12558_),
    .X(_12559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_694 ();
 sky130_fd_sc_hd__nor2_1 _18311_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(_12488_),
    .Y(_12561_));
 sky130_fd_sc_hd__a21oi_1 _18312_ (.A1(_12488_),
    .A2(_12559_),
    .B1(_12561_),
    .Y(_00279_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_693 ();
 sky130_fd_sc_hd__nor2_1 _18314_ (.A(_12285_),
    .B(_12435_),
    .Y(_12563_));
 sky130_fd_sc_hd__a211oi_1 _18315_ (.A1(\cs_registers_i.mstack_epc_q[2] ),
    .A2(_12400_),
    .B1(_12462_),
    .C1(_12563_),
    .Y(_12564_));
 sky130_fd_sc_hd__nor2_1 _18316_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .B(_12488_),
    .Y(_12565_));
 sky130_fd_sc_hd__a21oi_1 _18317_ (.A1(_12488_),
    .A2(_12564_),
    .B1(_12565_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _18318_ (.A(\cs_registers_i.mstack_epc_q[30] ),
    .B(_12400_),
    .Y(_12566_));
 sky130_fd_sc_hd__o221a_1 _18319_ (.A1(_12288_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11550_),
    .C1(_12566_),
    .X(_12567_));
 sky130_fd_sc_hd__nor2_1 _18320_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(_12488_),
    .Y(_12568_));
 sky130_fd_sc_hd__a21oi_1 _18321_ (.A1(_12488_),
    .A2(_12567_),
    .B1(_12568_),
    .Y(_00281_));
 sky130_fd_sc_hd__nor2_1 _18322_ (.A(_12291_),
    .B(_12435_),
    .Y(_12569_));
 sky130_fd_sc_hd__a211oi_1 _18323_ (.A1(\cs_registers_i.mstack_epc_q[31] ),
    .A2(_12400_),
    .B1(_12484_),
    .C1(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__nor2_1 _18324_ (.A(\cs_registers_i.csr_mepc_o[31] ),
    .B(_12488_),
    .Y(_12571_));
 sky130_fd_sc_hd__a21oi_1 _18325_ (.A1(_12488_),
    .A2(_12570_),
    .B1(_12571_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _18326_ (.A(\cs_registers_i.mstack_epc_q[3] ),
    .B(_12400_),
    .Y(_12572_));
 sky130_fd_sc_hd__o221a_1 _18327_ (.A1(_12294_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11612_),
    .C1(_12572_),
    .X(_12573_));
 sky130_fd_sc_hd__nor2_1 _18328_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(_12488_),
    .Y(_12574_));
 sky130_fd_sc_hd__a21oi_1 _18329_ (.A1(_12488_),
    .A2(_12573_),
    .B1(_12574_),
    .Y(_00283_));
 sky130_fd_sc_hd__nor2_1 _18330_ (.A(_12297_),
    .B(_12435_),
    .Y(_12575_));
 sky130_fd_sc_hd__a221oi_1 _18331_ (.A1(\cs_registers_i.mstack_epc_q[4] ),
    .A2(_12400_),
    .B1(_12402_),
    .B2(_11631_),
    .C1(_12575_),
    .Y(_12576_));
 sky130_fd_sc_hd__nor2_1 _18332_ (.A(\cs_registers_i.csr_mepc_o[4] ),
    .B(_12488_),
    .Y(_12577_));
 sky130_fd_sc_hd__a21oi_1 _18333_ (.A1(_12488_),
    .A2(_12576_),
    .B1(_12577_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _18334_ (.A(\cs_registers_i.mstack_epc_q[5] ),
    .B(_12400_),
    .Y(_12578_));
 sky130_fd_sc_hd__o221a_1 _18335_ (.A1(_12300_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11647_),
    .C1(_12578_),
    .X(_12579_));
 sky130_fd_sc_hd__nor2_1 _18336_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .B(_12488_),
    .Y(_12580_));
 sky130_fd_sc_hd__a21oi_1 _18337_ (.A1(_12488_),
    .A2(_12579_),
    .B1(_12580_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _18338_ (.A(\cs_registers_i.mstack_epc_q[6] ),
    .B(_12400_),
    .Y(_12581_));
 sky130_fd_sc_hd__o221a_1 _18339_ (.A1(_12303_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11664_),
    .C1(_12581_),
    .X(_12582_));
 sky130_fd_sc_hd__nor2_1 _18340_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(_12488_),
    .Y(_12583_));
 sky130_fd_sc_hd__a21oi_1 _18341_ (.A1(_12488_),
    .A2(_12582_),
    .B1(_12583_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _18342_ (.A(\cs_registers_i.mstack_epc_q[7] ),
    .B(_12400_),
    .Y(_12584_));
 sky130_fd_sc_hd__o221a_1 _18343_ (.A1(_12306_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11685_),
    .C1(_12584_),
    .X(_12585_));
 sky130_fd_sc_hd__nor2_1 _18344_ (.A(\cs_registers_i.csr_mepc_o[7] ),
    .B(_12488_),
    .Y(_12586_));
 sky130_fd_sc_hd__a21oi_1 _18345_ (.A1(_12488_),
    .A2(_12585_),
    .B1(_12586_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _18346_ (.A(\cs_registers_i.mstack_epc_q[8] ),
    .B(_12400_),
    .Y(_12587_));
 sky130_fd_sc_hd__o221a_1 _18347_ (.A1(_12309_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11707_),
    .C1(_12587_),
    .X(_12588_));
 sky130_fd_sc_hd__nor2_1 _18348_ (.A(\cs_registers_i.csr_mepc_o[8] ),
    .B(_12488_),
    .Y(_12589_));
 sky130_fd_sc_hd__a21oi_1 _18349_ (.A1(_12488_),
    .A2(_12588_),
    .B1(_12589_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _18350_ (.A(\cs_registers_i.mstack_epc_q[9] ),
    .B(_12400_),
    .Y(_12590_));
 sky130_fd_sc_hd__o221a_1 _18351_ (.A1(_12312_),
    .A2(_12435_),
    .B1(_12406_),
    .B2(_11726_),
    .C1(_12590_),
    .X(_12591_));
 sky130_fd_sc_hd__nor2_1 _18352_ (.A(\cs_registers_i.csr_mepc_o[9] ),
    .B(_12488_),
    .Y(_12592_));
 sky130_fd_sc_hd__a21oi_1 _18353_ (.A1(_12488_),
    .A2(_12591_),
    .B1(_12592_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_8 _18354_ (.A(_10620_),
    .B(net3501),
    .Y(_12593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_691 ();
 sky130_fd_sc_hd__nand2_1 _18357_ (.A(\cs_registers_i.mie_q[0] ),
    .B(_12593_),
    .Y(_12596_));
 sky130_fd_sc_hd__o21ai_0 _18358_ (.A1(_11270_),
    .A2(_12593_),
    .B1(_12596_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(\cs_registers_i.mie_q[10] ),
    .B(_12593_),
    .Y(_12597_));
 sky130_fd_sc_hd__o21ai_0 _18360_ (.A1(_11476_),
    .A2(_12593_),
    .B1(_12597_),
    .Y(_00291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_690 ();
 sky130_fd_sc_hd__nand2_1 _18362_ (.A(\cs_registers_i.mie_q[11] ),
    .B(_12593_),
    .Y(_12599_));
 sky130_fd_sc_hd__o21ai_0 _18363_ (.A1(_11490_),
    .A2(_12593_),
    .B1(_12599_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _18364_ (.A(\cs_registers_i.mie_q[12] ),
    .B(_12593_),
    .Y(_12600_));
 sky130_fd_sc_hd__o21ai_0 _18365_ (.A1(_11506_),
    .A2(_12593_),
    .B1(_12600_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _18366_ (.A(\cs_registers_i.mie_q[13] ),
    .B(_12593_),
    .Y(_12601_));
 sky130_fd_sc_hd__o21ai_0 _18367_ (.A1(_11530_),
    .A2(_12593_),
    .B1(_12601_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(\cs_registers_i.mie_q[14] ),
    .B(_12593_),
    .Y(_12602_));
 sky130_fd_sc_hd__o21ai_0 _18369_ (.A1(_11550_),
    .A2(_12593_),
    .B1(_12602_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(\cs_registers_i.mie_q[15] ),
    .B(_12593_),
    .Y(_12603_));
 sky130_fd_sc_hd__o21ai_0 _18371_ (.A1(_11177_),
    .A2(_12593_),
    .B1(_12603_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _18372_ (.A(\cs_registers_i.mie_q[16] ),
    .B(_12593_),
    .Y(_12604_));
 sky130_fd_sc_hd__o21ai_0 _18373_ (.A1(_11685_),
    .A2(_12593_),
    .B1(_12604_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _18374_ (.A(\cs_registers_i.mie_q[17] ),
    .B(_12593_),
    .Y(_12605_));
 sky130_fd_sc_hd__o21ai_0 _18375_ (.A1(_11612_),
    .A2(_12593_),
    .B1(_12605_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _18376_ (.A(\cs_registers_i.mie_q[1] ),
    .B(_12593_),
    .Y(_12606_));
 sky130_fd_sc_hd__o21ai_0 _18377_ (.A1(_11294_),
    .A2(_12593_),
    .B1(_12606_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _18378_ (.A(\cs_registers_i.mie_q[2] ),
    .B(_12593_),
    .Y(_12607_));
 sky130_fd_sc_hd__o21ai_0 _18379_ (.A1(_11319_),
    .A2(_12593_),
    .B1(_12607_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _18380_ (.A(\cs_registers_i.mie_q[3] ),
    .B(_12593_),
    .Y(_12608_));
 sky130_fd_sc_hd__o21ai_0 _18381_ (.A1(_11333_),
    .A2(_12593_),
    .B1(_12608_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(\cs_registers_i.mie_q[4] ),
    .B(_12593_),
    .Y(_12609_));
 sky130_fd_sc_hd__o21ai_0 _18383_ (.A1(_11369_),
    .A2(_12593_),
    .B1(_12609_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _18384_ (.A(\cs_registers_i.mie_q[5] ),
    .B(_12593_),
    .Y(_12610_));
 sky130_fd_sc_hd__o21ai_0 _18385_ (.A1(_11390_),
    .A2(_12593_),
    .B1(_12610_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(\cs_registers_i.mie_q[6] ),
    .B(_12593_),
    .Y(_12611_));
 sky130_fd_sc_hd__o21ai_0 _18387_ (.A1(_11406_),
    .A2(_12593_),
    .B1(_12611_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _18388_ (.A(\cs_registers_i.mie_q[7] ),
    .B(_12593_),
    .Y(_12612_));
 sky130_fd_sc_hd__o21ai_0 _18389_ (.A1(net3492),
    .A2(_12593_),
    .B1(_12612_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(\cs_registers_i.mie_q[8] ),
    .B(_12593_),
    .Y(_12613_));
 sky130_fd_sc_hd__o21ai_0 _18391_ (.A1(_11441_),
    .A2(_12593_),
    .B1(_12613_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _18392_ (.A(\cs_registers_i.mie_q[9] ),
    .B(_12593_),
    .Y(_12614_));
 sky130_fd_sc_hd__o21ai_0 _18393_ (.A1(_11457_),
    .A2(_12593_),
    .B1(_12614_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_8 _18394_ (.A(net3540),
    .B(net3501),
    .Y(_12615_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_688 ();
 sky130_fd_sc_hd__nand2_1 _18397_ (.A(\cs_registers_i.mscratch_q[0] ),
    .B(_12615_),
    .Y(_12618_));
 sky130_fd_sc_hd__o21ai_0 _18398_ (.A1(_11042_),
    .A2(_12615_),
    .B1(_12618_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _18399_ (.A(\cs_registers_i.mscratch_q[10] ),
    .B(_12615_),
    .Y(_12619_));
 sky130_fd_sc_hd__o21ai_0 _18400_ (.A1(_11145_),
    .A2(_12615_),
    .B1(_12619_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _18401_ (.A(\cs_registers_i.mscratch_q[11] ),
    .B(_12615_),
    .Y(_12620_));
 sky130_fd_sc_hd__o21ai_0 _18402_ (.A1(_11177_),
    .A2(_12615_),
    .B1(_12620_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _18403_ (.A(\cs_registers_i.mscratch_q[12] ),
    .B(_12615_),
    .Y(_12621_));
 sky130_fd_sc_hd__o21ai_0 _18404_ (.A1(_11197_),
    .A2(_12615_),
    .B1(_12621_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _18405_ (.A(\cs_registers_i.mscratch_q[13] ),
    .B(_12615_),
    .Y(_12622_));
 sky130_fd_sc_hd__o21ai_0 _18406_ (.A1(_11214_),
    .A2(_12615_),
    .B1(_12622_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _18407_ (.A(\cs_registers_i.mscratch_q[14] ),
    .B(_12615_),
    .Y(_12623_));
 sky130_fd_sc_hd__o21ai_0 _18408_ (.A1(_11235_),
    .A2(_12615_),
    .B1(_12623_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand2_1 _18409_ (.A(\cs_registers_i.mscratch_q[15] ),
    .B(_12615_),
    .Y(_12624_));
 sky130_fd_sc_hd__o21ai_0 _18410_ (.A1(_11255_),
    .A2(_12615_),
    .B1(_12624_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _18411_ (.A(\cs_registers_i.mscratch_q[16] ),
    .B(_12615_),
    .Y(_12625_));
 sky130_fd_sc_hd__o21ai_0 _18412_ (.A1(_11270_),
    .A2(_12615_),
    .B1(_12625_),
    .Y(_00315_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_687 ();
 sky130_fd_sc_hd__nand2_1 _18414_ (.A(\cs_registers_i.mscratch_q[17] ),
    .B(_12615_),
    .Y(_12627_));
 sky130_fd_sc_hd__o21ai_0 _18415_ (.A1(_11294_),
    .A2(_12615_),
    .B1(_12627_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _18416_ (.A(\cs_registers_i.mscratch_q[18] ),
    .B(_12615_),
    .Y(_12628_));
 sky130_fd_sc_hd__o21ai_0 _18417_ (.A1(_11319_),
    .A2(_12615_),
    .B1(_12628_),
    .Y(_00317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_686 ();
 sky130_fd_sc_hd__nand2_1 _18419_ (.A(\cs_registers_i.mscratch_q[19] ),
    .B(_12615_),
    .Y(_12630_));
 sky130_fd_sc_hd__o21ai_0 _18420_ (.A1(_11333_),
    .A2(_12615_),
    .B1(_12630_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _18421_ (.A(\cs_registers_i.mscratch_q[1] ),
    .B(_12615_),
    .Y(_12631_));
 sky130_fd_sc_hd__o21ai_0 _18422_ (.A1(_11354_),
    .A2(_12615_),
    .B1(_12631_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _18423_ (.A(\cs_registers_i.mscratch_q[20] ),
    .B(_12615_),
    .Y(_12632_));
 sky130_fd_sc_hd__o21ai_0 _18424_ (.A1(_11369_),
    .A2(_12615_),
    .B1(_12632_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _18425_ (.A(\cs_registers_i.mscratch_q[21] ),
    .B(_12615_),
    .Y(_12633_));
 sky130_fd_sc_hd__o21ai_0 _18426_ (.A1(_11390_),
    .A2(_12615_),
    .B1(_12633_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(\cs_registers_i.mscratch_q[22] ),
    .B(_12615_),
    .Y(_12634_));
 sky130_fd_sc_hd__o21ai_0 _18428_ (.A1(_11406_),
    .A2(_12615_),
    .B1(_12634_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _18429_ (.A(\cs_registers_i.mscratch_q[23] ),
    .B(_12615_),
    .Y(_12635_));
 sky130_fd_sc_hd__o21ai_0 _18430_ (.A1(_11426_),
    .A2(_12615_),
    .B1(_12635_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(\cs_registers_i.mscratch_q[24] ),
    .B(_12615_),
    .Y(_12636_));
 sky130_fd_sc_hd__o21ai_0 _18432_ (.A1(_11441_),
    .A2(_12615_),
    .B1(_12636_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _18433_ (.A(\cs_registers_i.mscratch_q[25] ),
    .B(_12615_),
    .Y(_12637_));
 sky130_fd_sc_hd__o21ai_0 _18434_ (.A1(_11457_),
    .A2(_12615_),
    .B1(_12637_),
    .Y(_00325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_685 ();
 sky130_fd_sc_hd__nand2_1 _18436_ (.A(\cs_registers_i.mscratch_q[26] ),
    .B(_12615_),
    .Y(_12639_));
 sky130_fd_sc_hd__o21ai_0 _18437_ (.A1(_11476_),
    .A2(_12615_),
    .B1(_12639_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _18438_ (.A(\cs_registers_i.mscratch_q[27] ),
    .B(_12615_),
    .Y(_12640_));
 sky130_fd_sc_hd__o21ai_0 _18439_ (.A1(_11490_),
    .A2(_12615_),
    .B1(_12640_),
    .Y(_00327_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_684 ();
 sky130_fd_sc_hd__nand2_1 _18441_ (.A(\cs_registers_i.mscratch_q[28] ),
    .B(_12615_),
    .Y(_12642_));
 sky130_fd_sc_hd__o21ai_0 _18442_ (.A1(_11506_),
    .A2(_12615_),
    .B1(_12642_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _18443_ (.A(\cs_registers_i.mscratch_q[29] ),
    .B(_12615_),
    .Y(_12643_));
 sky130_fd_sc_hd__o21ai_0 _18444_ (.A1(_11530_),
    .A2(_12615_),
    .B1(_12643_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _18445_ (.A(\cs_registers_i.mscratch_q[2] ),
    .B(_12615_),
    .Y(_12644_));
 sky130_fd_sc_hd__o21ai_0 _18446_ (.A1(_11082_),
    .A2(_12615_),
    .B1(_12644_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _18447_ (.A(\cs_registers_i.mscratch_q[30] ),
    .B(_12615_),
    .Y(_12645_));
 sky130_fd_sc_hd__o21ai_0 _18448_ (.A1(_11550_),
    .A2(_12615_),
    .B1(_12645_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _18449_ (.A(\cs_registers_i.mscratch_q[31] ),
    .B(_12615_),
    .Y(_12646_));
 sky130_fd_sc_hd__o21ai_0 _18450_ (.A1(_11565_),
    .A2(_12615_),
    .B1(_12646_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _18451_ (.A(\cs_registers_i.mscratch_q[3] ),
    .B(_12615_),
    .Y(_12647_));
 sky130_fd_sc_hd__o21ai_0 _18452_ (.A1(_11612_),
    .A2(_12615_),
    .B1(_12647_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(\cs_registers_i.mscratch_q[4] ),
    .B(_12615_),
    .Y(_12648_));
 sky130_fd_sc_hd__o21ai_0 _18454_ (.A1(_11780_),
    .A2(_12615_),
    .B1(_12648_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _18455_ (.A(\cs_registers_i.mscratch_q[5] ),
    .B(_12615_),
    .Y(_12649_));
 sky130_fd_sc_hd__o21ai_0 _18456_ (.A1(_11647_),
    .A2(_12615_),
    .B1(_12649_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _18457_ (.A(\cs_registers_i.mscratch_q[6] ),
    .B(_12615_),
    .Y(_12650_));
 sky130_fd_sc_hd__o21ai_0 _18458_ (.A1(_11664_),
    .A2(_12615_),
    .B1(_12650_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _18459_ (.A(\cs_registers_i.mscratch_q[7] ),
    .B(_12615_),
    .Y(_12651_));
 sky130_fd_sc_hd__o21ai_0 _18460_ (.A1(net3478),
    .A2(_12615_),
    .B1(_12651_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _18461_ (.A(\cs_registers_i.mscratch_q[8] ),
    .B(_12615_),
    .Y(_12652_));
 sky130_fd_sc_hd__o21ai_0 _18462_ (.A1(_11707_),
    .A2(_12615_),
    .B1(_12652_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(\cs_registers_i.mscratch_q[9] ),
    .B(_12615_),
    .Y(_12653_));
 sky130_fd_sc_hd__o21ai_0 _18464_ (.A1(_11726_),
    .A2(_12615_),
    .B1(_12653_),
    .Y(_00339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_683 ();
 sky130_fd_sc_hd__nand2_1 _18466_ (.A(\cs_registers_i.mcause_q[0] ),
    .B(net3532),
    .Y(_12655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_682 ();
 sky130_fd_sc_hd__nand2_1 _18468_ (.A(\cs_registers_i.mstack_cause_q[0] ),
    .B(_12435_),
    .Y(_12657_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(_12655_),
    .B(_12657_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _18470_ (.A(\cs_registers_i.mcause_q[1] ),
    .B(_12394_),
    .Y(_12658_));
 sky130_fd_sc_hd__nand2_1 _18471_ (.A(\cs_registers_i.mstack_cause_q[1] ),
    .B(_12435_),
    .Y(_12659_));
 sky130_fd_sc_hd__nand2_1 _18472_ (.A(_12658_),
    .B(_12659_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _18473_ (.A(\cs_registers_i.mcause_q[2] ),
    .B(_12394_),
    .Y(_12660_));
 sky130_fd_sc_hd__nand2_1 _18474_ (.A(\cs_registers_i.mstack_cause_q[2] ),
    .B(_12435_),
    .Y(_12661_));
 sky130_fd_sc_hd__nand2_1 _18475_ (.A(_12660_),
    .B(_12661_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _18476_ (.A(\cs_registers_i.mcause_q[3] ),
    .B(net3532),
    .Y(_12662_));
 sky130_fd_sc_hd__nand2_1 _18477_ (.A(\cs_registers_i.mstack_cause_q[3] ),
    .B(_12435_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_1 _18478_ (.A(_12662_),
    .B(_12663_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _18479_ (.A(\cs_registers_i.mcause_q[4] ),
    .B(net3532),
    .Y(_12664_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(\cs_registers_i.mstack_cause_q[4] ),
    .B(_12435_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand2_1 _18481_ (.A(_12664_),
    .B(_12665_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(\cs_registers_i.mcause_q[5] ),
    .B(_12394_),
    .Y(_12666_));
 sky130_fd_sc_hd__nand2_1 _18483_ (.A(\cs_registers_i.mstack_cause_q[5] ),
    .B(_12435_),
    .Y(_12667_));
 sky130_fd_sc_hd__nand2_1 _18484_ (.A(_12666_),
    .B(_12667_),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _18485_ (.A(\cs_registers_i.mstatus_q[2] ),
    .B(net3532),
    .Y(_12668_));
 sky130_fd_sc_hd__nand2_1 _18486_ (.A(\cs_registers_i.mstack_q[0] ),
    .B(_12435_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_12668_),
    .B(_12669_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(\cs_registers_i.mstatus_q[3] ),
    .B(_12394_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(\cs_registers_i.mstack_q[1] ),
    .B(_12435_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_1 _18490_ (.A(_12670_),
    .B(_12671_),
    .Y(_00347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_680 ();
 sky130_fd_sc_hd__nand2_1 _18493_ (.A(\cs_registers_i.mstatus_q[4] ),
    .B(net3532),
    .Y(_12674_));
 sky130_fd_sc_hd__nand2_1 _18494_ (.A(\cs_registers_i.mstack_q[2] ),
    .B(_12435_),
    .Y(_12675_));
 sky130_fd_sc_hd__nand2_1 _18495_ (.A(_12674_),
    .B(_12675_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _18496_ (.A(\cs_registers_i.csr_mepc_o[0] ),
    .B(net3532),
    .Y(_12676_));
 sky130_fd_sc_hd__nand2_1 _18497_ (.A(\cs_registers_i.mstack_epc_q[0] ),
    .B(_12435_),
    .Y(_12677_));
 sky130_fd_sc_hd__nand2_1 _18498_ (.A(_12676_),
    .B(_12677_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _18499_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(_12394_),
    .Y(_12678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_679 ();
 sky130_fd_sc_hd__nand2_1 _18501_ (.A(\cs_registers_i.mstack_epc_q[10] ),
    .B(_12435_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand2_1 _18502_ (.A(_12678_),
    .B(_12680_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _18503_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(net3532),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_1 _18504_ (.A(\cs_registers_i.mstack_epc_q[11] ),
    .B(_12435_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand2_1 _18505_ (.A(_12681_),
    .B(_12682_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _18506_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(_12394_),
    .Y(_12683_));
 sky130_fd_sc_hd__nand2_1 _18507_ (.A(\cs_registers_i.mstack_epc_q[12] ),
    .B(_12435_),
    .Y(_12684_));
 sky130_fd_sc_hd__nand2_1 _18508_ (.A(_12683_),
    .B(_12684_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _18509_ (.A(\cs_registers_i.csr_mepc_o[13] ),
    .B(_12394_),
    .Y(_12685_));
 sky130_fd_sc_hd__nand2_1 _18510_ (.A(\cs_registers_i.mstack_epc_q[13] ),
    .B(_12435_),
    .Y(_12686_));
 sky130_fd_sc_hd__nand2_1 _18511_ (.A(_12685_),
    .B(_12686_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _18512_ (.A(\cs_registers_i.csr_mepc_o[14] ),
    .B(net3532),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_1 _18513_ (.A(\cs_registers_i.mstack_epc_q[14] ),
    .B(_12435_),
    .Y(_12688_));
 sky130_fd_sc_hd__nand2_1 _18514_ (.A(_12687_),
    .B(_12688_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _18515_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(_12394_),
    .Y(_12689_));
 sky130_fd_sc_hd__nand2_1 _18516_ (.A(\cs_registers_i.mstack_epc_q[15] ),
    .B(_12435_),
    .Y(_12690_));
 sky130_fd_sc_hd__nand2_1 _18517_ (.A(_12689_),
    .B(_12690_),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _18518_ (.A(\cs_registers_i.csr_mepc_o[16] ),
    .B(_12394_),
    .Y(_12691_));
 sky130_fd_sc_hd__nand2_1 _18519_ (.A(\cs_registers_i.mstack_epc_q[16] ),
    .B(_12435_),
    .Y(_12692_));
 sky130_fd_sc_hd__nand2_1 _18520_ (.A(_12691_),
    .B(_12692_),
    .Y(_00356_));
 sky130_fd_sc_hd__nand2_1 _18521_ (.A(\cs_registers_i.csr_mepc_o[17] ),
    .B(_12394_),
    .Y(_12693_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(\cs_registers_i.mstack_epc_q[17] ),
    .B(_12435_),
    .Y(_12694_));
 sky130_fd_sc_hd__nand2_1 _18523_ (.A(_12693_),
    .B(_12694_),
    .Y(_00357_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_678 ();
 sky130_fd_sc_hd__nand2_1 _18525_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(net3532),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_1 _18526_ (.A(\cs_registers_i.mstack_epc_q[18] ),
    .B(_12435_),
    .Y(_12697_));
 sky130_fd_sc_hd__nand2_1 _18527_ (.A(_12696_),
    .B(_12697_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2_1 _18528_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(net3532),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_1 _18529_ (.A(\cs_registers_i.mstack_epc_q[19] ),
    .B(_12435_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand2_1 _18530_ (.A(_12698_),
    .B(_12699_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _18531_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(_12394_),
    .Y(_12700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_677 ();
 sky130_fd_sc_hd__nand2_1 _18533_ (.A(\cs_registers_i.mstack_epc_q[1] ),
    .B(_12435_),
    .Y(_12702_));
 sky130_fd_sc_hd__nand2_1 _18534_ (.A(_12700_),
    .B(_12702_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _18535_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(net3532),
    .Y(_12703_));
 sky130_fd_sc_hd__nand2_1 _18536_ (.A(\cs_registers_i.mstack_epc_q[20] ),
    .B(_12435_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand2_1 _18537_ (.A(_12703_),
    .B(_12704_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _18538_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(net3532),
    .Y(_12705_));
 sky130_fd_sc_hd__nand2_1 _18539_ (.A(\cs_registers_i.mstack_epc_q[21] ),
    .B(_12435_),
    .Y(_12706_));
 sky130_fd_sc_hd__nand2_1 _18540_ (.A(_12705_),
    .B(_12706_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _18541_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(net3532),
    .Y(_12707_));
 sky130_fd_sc_hd__nand2_1 _18542_ (.A(\cs_registers_i.mstack_epc_q[22] ),
    .B(_12435_),
    .Y(_12708_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(_12707_),
    .B(_12708_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _18544_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(net3532),
    .Y(_12709_));
 sky130_fd_sc_hd__nand2_1 _18545_ (.A(\cs_registers_i.mstack_epc_q[23] ),
    .B(_12435_),
    .Y(_12710_));
 sky130_fd_sc_hd__nand2_1 _18546_ (.A(_12709_),
    .B(_12710_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(net3532),
    .Y(_12711_));
 sky130_fd_sc_hd__nand2_1 _18548_ (.A(\cs_registers_i.mstack_epc_q[24] ),
    .B(_12435_),
    .Y(_12712_));
 sky130_fd_sc_hd__nand2_1 _18549_ (.A(_12711_),
    .B(_12712_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _18550_ (.A(\cs_registers_i.csr_mepc_o[25] ),
    .B(net3532),
    .Y(_12713_));
 sky130_fd_sc_hd__nand2_1 _18551_ (.A(\cs_registers_i.mstack_epc_q[25] ),
    .B(_12435_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(_12713_),
    .B(_12714_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _18553_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(net3532),
    .Y(_12715_));
 sky130_fd_sc_hd__nand2_1 _18554_ (.A(\cs_registers_i.mstack_epc_q[26] ),
    .B(_12435_),
    .Y(_12716_));
 sky130_fd_sc_hd__nand2_1 _18555_ (.A(_12715_),
    .B(_12716_),
    .Y(_00367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_676 ();
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(net3532),
    .Y(_12718_));
 sky130_fd_sc_hd__nand2_1 _18558_ (.A(\cs_registers_i.mstack_epc_q[27] ),
    .B(_12435_),
    .Y(_12719_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(_12718_),
    .B(_12719_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(\cs_registers_i.csr_mepc_o[28] ),
    .B(net3532),
    .Y(_12720_));
 sky130_fd_sc_hd__nand2_1 _18561_ (.A(\cs_registers_i.mstack_epc_q[28] ),
    .B(_12435_),
    .Y(_12721_));
 sky130_fd_sc_hd__nand2_1 _18562_ (.A(_12720_),
    .B(_12721_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _18563_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(net3532),
    .Y(_12722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_675 ();
 sky130_fd_sc_hd__nand2_1 _18565_ (.A(\cs_registers_i.mstack_epc_q[29] ),
    .B(_12435_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand2_1 _18566_ (.A(_12722_),
    .B(_12724_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(\cs_registers_i.mstack_epc_q[2] ),
    .B(_12435_),
    .Y(_12725_));
 sky130_fd_sc_hd__o21ai_0 _18568_ (.A1(_11073_),
    .A2(_12435_),
    .B1(_12725_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(net3532),
    .Y(_12726_));
 sky130_fd_sc_hd__nand2_1 _18570_ (.A(\cs_registers_i.mstack_epc_q[30] ),
    .B(_12435_),
    .Y(_12727_));
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(_12726_),
    .B(_12727_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_1 _18572_ (.A(\cs_registers_i.csr_mepc_o[31] ),
    .B(_12394_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand2_1 _18573_ (.A(\cs_registers_i.mstack_epc_q[31] ),
    .B(_12435_),
    .Y(_12729_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(_12728_),
    .B(_12729_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _18575_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(net3532),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_1 _18576_ (.A(\cs_registers_i.mstack_epc_q[3] ),
    .B(_12435_),
    .Y(_12731_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(_12730_),
    .B(_12731_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(\cs_registers_i.csr_mepc_o[4] ),
    .B(_12394_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand2_1 _18579_ (.A(\cs_registers_i.mstack_epc_q[4] ),
    .B(_12435_),
    .Y(_12733_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(_12732_),
    .B(_12733_),
    .Y(_00375_));
 sky130_fd_sc_hd__nand2_1 _18581_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .B(_12394_),
    .Y(_12734_));
 sky130_fd_sc_hd__nand2_1 _18582_ (.A(\cs_registers_i.mstack_epc_q[5] ),
    .B(_12435_),
    .Y(_12735_));
 sky130_fd_sc_hd__nand2_1 _18583_ (.A(_12734_),
    .B(_12735_),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(_12394_),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_1 _18585_ (.A(\cs_registers_i.mstack_epc_q[6] ),
    .B(_12435_),
    .Y(_12737_));
 sky130_fd_sc_hd__nand2_1 _18586_ (.A(_12736_),
    .B(_12737_),
    .Y(_00377_));
 sky130_fd_sc_hd__nand2_1 _18587_ (.A(\cs_registers_i.csr_mepc_o[7] ),
    .B(_12394_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(\cs_registers_i.mstack_epc_q[7] ),
    .B(_12435_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(_12738_),
    .B(_12739_),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _18590_ (.A(\cs_registers_i.csr_mepc_o[8] ),
    .B(_12394_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_1 _18591_ (.A(\cs_registers_i.mstack_epc_q[8] ),
    .B(_12435_),
    .Y(_12741_));
 sky130_fd_sc_hd__nand2_1 _18592_ (.A(_12740_),
    .B(_12741_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _18593_ (.A(\cs_registers_i.csr_mepc_o[9] ),
    .B(_12394_),
    .Y(_12742_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(\cs_registers_i.mstack_epc_q[9] ),
    .B(_12435_),
    .Y(_12743_));
 sky130_fd_sc_hd__nand2_1 _18595_ (.A(_12742_),
    .B(_12743_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2_2 _18596_ (.A(_10595_),
    .B(net3501),
    .Y(_12744_));
 sky130_fd_sc_hd__nand2_1 _18597_ (.A(\cs_registers_i.csr_mstatus_tw_o ),
    .B(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__o21ai_0 _18598_ (.A1(_11390_),
    .A2(_12744_),
    .B1(_12745_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(\cs_registers_i.mstatus_q[1] ),
    .B(_12744_),
    .Y(_12746_));
 sky130_fd_sc_hd__o21ai_0 _18600_ (.A1(_11294_),
    .A2(_12744_),
    .B1(_12746_),
    .Y(_00382_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_674 ();
 sky130_fd_sc_hd__nand2_8 _18602_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_10646_),
    .Y(_12748_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_672 ();
 sky130_fd_sc_hd__mux2i_1 _18605_ (.A0(net329),
    .A1(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(net3947),
    .Y(_12751_));
 sky130_fd_sc_hd__nor2_1 _18606_ (.A(_12748_),
    .B(_12751_),
    .Y(_12752_));
 sky130_fd_sc_hd__a21oi_1 _18607_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(net3609),
    .B1(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__and3_4 _18608_ (.A(_10495_),
    .B(_10499_),
    .C(_10784_),
    .X(_12754_));
 sky130_fd_sc_hd__o311ai_1 _18609_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_12416_),
    .A3(net3609),
    .B1(_12394_),
    .C1(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_671 ();
 sky130_fd_sc_hd__nand2_8 _18611_ (.A(net3539),
    .B(net3501),
    .Y(_12757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_669 ();
 sky130_fd_sc_hd__nor2_1 _18614_ (.A(_11042_),
    .B(_12757_),
    .Y(_12760_));
 sky130_fd_sc_hd__a21oi_1 _18615_ (.A1(\cs_registers_i.mtval_q[0] ),
    .A2(_12757_),
    .B1(_12760_),
    .Y(_12761_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_668 ();
 sky130_fd_sc_hd__o22ai_1 _18617_ (.A1(_12753_),
    .A2(net3524),
    .B1(_12761_),
    .B2(_12394_),
    .Y(_00387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_667 ();
 sky130_fd_sc_hd__mux2_8 _18619_ (.A0(net3946),
    .A1(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .S(net3947),
    .X(_12764_));
 sky130_fd_sc_hd__nand2_2 _18620_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Y(_12765_));
 sky130_fd_sc_hd__nor3_2 _18621_ (.A(_08414_),
    .B(_08404_),
    .C(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__and3_4 _18622_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(\cs_registers_i.pc_id_i[5] ),
    .C(_12766_),
    .X(_12767_));
 sky130_fd_sc_hd__and3_4 _18623_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(\cs_registers_i.pc_id_i[7] ),
    .C(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__nand3_2 _18624_ (.A(net3823),
    .B(\cs_registers_i.pc_id_i[9] ),
    .C(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__xnor2_1 _18625_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(_12769_),
    .Y(_12770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_666 ();
 sky130_fd_sc_hd__a222oi_1 _18627_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12764_),
    .C1(_12770_),
    .C2(_12416_),
    .Y(_12772_));
 sky130_fd_sc_hd__nor2_1 _18628_ (.A(_11145_),
    .B(_12757_),
    .Y(_12773_));
 sky130_fd_sc_hd__a21oi_1 _18629_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(_12757_),
    .B1(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__o22ai_1 _18630_ (.A1(net3524),
    .A2(_12772_),
    .B1(_12774_),
    .B2(_12394_),
    .Y(_00388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_664 ();
 sky130_fd_sc_hd__mux2_8 _18633_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .S(net3947),
    .X(_12777_));
 sky130_fd_sc_hd__inv_1 _18634_ (.A(\cs_registers_i.pc_id_i[10] ),
    .Y(_12778_));
 sky130_fd_sc_hd__nor2_2 _18635_ (.A(_12778_),
    .B(_12769_),
    .Y(_12779_));
 sky130_fd_sc_hd__xor2_1 _18636_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_12779_),
    .X(_12780_));
 sky130_fd_sc_hd__a222oi_1 _18637_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12777_),
    .C1(_12780_),
    .C2(_12416_),
    .Y(_12781_));
 sky130_fd_sc_hd__nor2_1 _18638_ (.A(_11177_),
    .B(_12757_),
    .Y(_12782_));
 sky130_fd_sc_hd__a21oi_1 _18639_ (.A1(\cs_registers_i.mtval_q[11] ),
    .A2(_12757_),
    .B1(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__o22ai_1 _18640_ (.A1(net3524),
    .A2(_12781_),
    .B1(_12783_),
    .B2(_12394_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(net3947),
    .B(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .Y(_12784_));
 sky130_fd_sc_hd__o21ai_0 _18642_ (.A1(_08008_),
    .A2(net3947),
    .B1(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_12779_),
    .Y(_12786_));
 sky130_fd_sc_hd__xnor2_1 _18644_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__a222oi_1 _18645_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12785_),
    .C1(_12787_),
    .C2(_12416_),
    .Y(_12788_));
 sky130_fd_sc_hd__nor2_1 _18646_ (.A(_11197_),
    .B(_12757_),
    .Y(_12789_));
 sky130_fd_sc_hd__a21oi_1 _18647_ (.A1(\cs_registers_i.mtval_q[12] ),
    .A2(_12757_),
    .B1(_12789_),
    .Y(_12790_));
 sky130_fd_sc_hd__o22ai_1 _18648_ (.A1(net3524),
    .A2(_12788_),
    .B1(_12790_),
    .B2(_12394_),
    .Y(_00390_));
 sky130_fd_sc_hd__mux2_4 _18649_ (.A0(net3938),
    .A1(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .S(net3947),
    .X(_12791_));
 sky130_fd_sc_hd__nand3_2 _18650_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(\cs_registers_i.pc_id_i[11] ),
    .C(_12779_),
    .Y(_12792_));
 sky130_fd_sc_hd__xnor2_1 _18651_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__a222oi_1 _18652_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12791_),
    .C1(_12793_),
    .C2(_12416_),
    .Y(_12794_));
 sky130_fd_sc_hd__nor2_1 _18653_ (.A(_11214_),
    .B(_12757_),
    .Y(_12795_));
 sky130_fd_sc_hd__a21oi_1 _18654_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(_12757_),
    .B1(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__o22ai_1 _18655_ (.A1(net3524),
    .A2(_12794_),
    .B1(_12796_),
    .B2(_12394_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_2 _18656_ (.A(net3947),
    .B(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .Y(_12797_));
 sky130_fd_sc_hd__o21ai_0 _18657_ (.A1(_08009_),
    .A2(net3947),
    .B1(_12797_),
    .Y(_12798_));
 sky130_fd_sc_hd__inv_1 _18658_ (.A(\cs_registers_i.pc_id_i[13] ),
    .Y(_12799_));
 sky130_fd_sc_hd__nor2_2 _18659_ (.A(_12799_),
    .B(_12792_),
    .Y(_12800_));
 sky130_fd_sc_hd__xor2_1 _18660_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(_12800_),
    .X(_12801_));
 sky130_fd_sc_hd__a222oi_1 _18661_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12798_),
    .C1(_12801_),
    .C2(_12416_),
    .Y(_12802_));
 sky130_fd_sc_hd__nor2_1 _18662_ (.A(_11235_),
    .B(_12757_),
    .Y(_12803_));
 sky130_fd_sc_hd__a21oi_1 _18663_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(_12757_),
    .B1(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__o22ai_1 _18664_ (.A1(net3524),
    .A2(_12802_),
    .B1(_12804_),
    .B2(net3532),
    .Y(_00392_));
 sky130_fd_sc_hd__mux2_8 _18665_ (.A0(net3933),
    .A1(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .S(net3947),
    .X(_12805_));
 sky130_fd_sc_hd__nand2_1 _18666_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(_12800_),
    .Y(_12806_));
 sky130_fd_sc_hd__xnor2_1 _18667_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_12806_),
    .Y(_12807_));
 sky130_fd_sc_hd__a222oi_1 _18668_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12805_),
    .C1(_12807_),
    .C2(_12416_),
    .Y(_12808_));
 sky130_fd_sc_hd__nor2_1 _18669_ (.A(_11255_),
    .B(_12757_),
    .Y(_12809_));
 sky130_fd_sc_hd__a21oi_1 _18670_ (.A1(\cs_registers_i.mtval_q[15] ),
    .A2(_12757_),
    .B1(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__o22ai_1 _18671_ (.A1(net3524),
    .A2(_12808_),
    .B1(_12810_),
    .B2(_12394_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand3_2 _18672_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(\cs_registers_i.pc_id_i[15] ),
    .C(_12800_),
    .Y(_12811_));
 sky130_fd_sc_hd__xnor2_1 _18673_ (.A(\cs_registers_i.pc_id_i[16] ),
    .B(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__nor2_4 _18674_ (.A(net3947),
    .B(_12748_),
    .Y(_12813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_663 ();
 sky130_fd_sc_hd__a222oi_1 _18676_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net3609),
    .B1(_12812_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3915),
    .Y(_12815_));
 sky130_fd_sc_hd__nor2_1 _18677_ (.A(_11270_),
    .B(_12757_),
    .Y(_12816_));
 sky130_fd_sc_hd__a21oi_1 _18678_ (.A1(\cs_registers_i.mtval_q[16] ),
    .A2(_12757_),
    .B1(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__o22ai_1 _18679_ (.A1(net3524),
    .A2(_12815_),
    .B1(_12817_),
    .B2(_12394_),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_1 _18680_ (.A(\cs_registers_i.pc_id_i[16] ),
    .Y(_12818_));
 sky130_fd_sc_hd__nor2_2 _18681_ (.A(_12818_),
    .B(_12811_),
    .Y(_12819_));
 sky130_fd_sc_hd__xor2_1 _18682_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_12819_),
    .X(_12820_));
 sky130_fd_sc_hd__a222oi_1 _18683_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net3609),
    .B1(_12820_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3901),
    .Y(_12821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_662 ();
 sky130_fd_sc_hd__nor2_1 _18685_ (.A(_11294_),
    .B(_12757_),
    .Y(_12823_));
 sky130_fd_sc_hd__a21oi_1 _18686_ (.A1(\cs_registers_i.mtval_q[17] ),
    .A2(_12757_),
    .B1(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__o22ai_1 _18687_ (.A1(net3524),
    .A2(_12821_),
    .B1(_12824_),
    .B2(_12394_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_12819_),
    .Y(_12825_));
 sky130_fd_sc_hd__xnor2_1 _18689_ (.A(\cs_registers_i.pc_id_i[18] ),
    .B(_12825_),
    .Y(_12826_));
 sky130_fd_sc_hd__a222oi_1 _18690_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net3609),
    .B1(_12826_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3897),
    .Y(_12827_));
 sky130_fd_sc_hd__nor2_1 _18691_ (.A(_11319_),
    .B(_12757_),
    .Y(_12828_));
 sky130_fd_sc_hd__a21oi_1 _18692_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_12757_),
    .B1(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__o22ai_1 _18693_ (.A1(net3524),
    .A2(_12827_),
    .B1(_12829_),
    .B2(net3532),
    .Y(_00396_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_661 ();
 sky130_fd_sc_hd__nand3_2 _18695_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(\cs_registers_i.pc_id_i[18] ),
    .C(_12819_),
    .Y(_12831_));
 sky130_fd_sc_hd__xnor2_1 _18696_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_660 ();
 sky130_fd_sc_hd__a222oi_1 _18698_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net3609),
    .B1(_12832_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3896),
    .Y(_12834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_659 ();
 sky130_fd_sc_hd__nor2_1 _18700_ (.A(_11333_),
    .B(_12757_),
    .Y(_12836_));
 sky130_fd_sc_hd__a21oi_1 _18701_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_12757_),
    .B1(_12836_),
    .Y(_12837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_658 ();
 sky130_fd_sc_hd__o22ai_1 _18703_ (.A1(net3524),
    .A2(_12834_),
    .B1(_12837_),
    .B2(_12394_),
    .Y(_00397_));
 sky130_fd_sc_hd__mux2i_1 _18704_ (.A0(\id_stage_i.controller_i.instr_i[1] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .S(net3947),
    .Y(_12839_));
 sky130_fd_sc_hd__xnor2_1 _18705_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Y(_12840_));
 sky130_fd_sc_hd__o22ai_1 _18706_ (.A1(_12748_),
    .A2(_12839_),
    .B1(_12840_),
    .B2(_10646_),
    .Y(_12841_));
 sky130_fd_sc_hd__a21oi_2 _18707_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(net3609),
    .B1(_12841_),
    .Y(_12842_));
 sky130_fd_sc_hd__nor2_1 _18708_ (.A(_11354_),
    .B(_12757_),
    .Y(_12843_));
 sky130_fd_sc_hd__a21oi_1 _18709_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(_12757_),
    .B1(_12843_),
    .Y(_12844_));
 sky130_fd_sc_hd__o22ai_1 _18710_ (.A1(net3524),
    .A2(_12842_),
    .B1(_12844_),
    .B2(_12394_),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_1 _18711_ (.A(\cs_registers_i.pc_id_i[19] ),
    .Y(_12845_));
 sky130_fd_sc_hd__nor2_2 _18712_ (.A(_12845_),
    .B(_12831_),
    .Y(_12846_));
 sky130_fd_sc_hd__xor2_1 _18713_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(_12846_),
    .X(_12847_));
 sky130_fd_sc_hd__a222oi_1 _18714_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net3609),
    .B1(_12847_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3895),
    .Y(_12848_));
 sky130_fd_sc_hd__nor2_1 _18715_ (.A(_11369_),
    .B(_12757_),
    .Y(_12849_));
 sky130_fd_sc_hd__a21oi_1 _18716_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_12757_),
    .B1(_12849_),
    .Y(_12850_));
 sky130_fd_sc_hd__o22ai_1 _18717_ (.A1(net3524),
    .A2(_12848_),
    .B1(_12850_),
    .B2(net3532),
    .Y(_00399_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_657 ();
 sky130_fd_sc_hd__nand2_1 _18719_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(_12846_),
    .Y(_12852_));
 sky130_fd_sc_hd__xnor2_1 _18720_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(_12852_),
    .Y(_12853_));
 sky130_fd_sc_hd__a222oi_1 _18721_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net3609),
    .B1(_12853_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3858),
    .Y(_12854_));
 sky130_fd_sc_hd__nor2_1 _18722_ (.A(_11390_),
    .B(_12757_),
    .Y(_12855_));
 sky130_fd_sc_hd__a21oi_1 _18723_ (.A1(\cs_registers_i.mtval_q[21] ),
    .A2(_12757_),
    .B1(_12855_),
    .Y(_12856_));
 sky130_fd_sc_hd__o22ai_1 _18724_ (.A1(net3524),
    .A2(_12854_),
    .B1(_12856_),
    .B2(_12394_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand3_2 _18725_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(\cs_registers_i.pc_id_i[21] ),
    .C(_12846_),
    .Y(_12857_));
 sky130_fd_sc_hd__xnor2_1 _18726_ (.A(\cs_registers_i.pc_id_i[22] ),
    .B(_12857_),
    .Y(_12858_));
 sky130_fd_sc_hd__a222oi_1 _18727_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net3609),
    .B1(_12858_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3851),
    .Y(_12859_));
 sky130_fd_sc_hd__nor2_1 _18728_ (.A(_11406_),
    .B(_12757_),
    .Y(_12860_));
 sky130_fd_sc_hd__a21oi_1 _18729_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_12757_),
    .B1(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__o22ai_1 _18730_ (.A1(net3524),
    .A2(_12859_),
    .B1(_12861_),
    .B2(_12394_),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_1 _18731_ (.A(\cs_registers_i.pc_id_i[22] ),
    .Y(_12862_));
 sky130_fd_sc_hd__nor2_2 _18732_ (.A(_12862_),
    .B(_12857_),
    .Y(_12863_));
 sky130_fd_sc_hd__xor2_1 _18733_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_12863_),
    .X(_12864_));
 sky130_fd_sc_hd__a222oi_1 _18734_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net3609),
    .B1(_12864_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net285),
    .Y(_12865_));
 sky130_fd_sc_hd__nor2_1 _18735_ (.A(_11426_),
    .B(_12757_),
    .Y(_12866_));
 sky130_fd_sc_hd__a21oi_1 _18736_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_12757_),
    .B1(_12866_),
    .Y(_12867_));
 sky130_fd_sc_hd__o22ai_1 _18737_ (.A1(net3524),
    .A2(_12865_),
    .B1(_12867_),
    .B2(_12394_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _18738_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_12863_),
    .Y(_12868_));
 sky130_fd_sc_hd__xnor2_1 _18739_ (.A(\cs_registers_i.pc_id_i[24] ),
    .B(_12868_),
    .Y(_12869_));
 sky130_fd_sc_hd__a222oi_1 _18740_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net3609),
    .B1(_12869_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3845),
    .Y(_12870_));
 sky130_fd_sc_hd__nor2_1 _18741_ (.A(_11441_),
    .B(_12757_),
    .Y(_12871_));
 sky130_fd_sc_hd__a21oi_1 _18742_ (.A1(\cs_registers_i.mtval_q[24] ),
    .A2(_12757_),
    .B1(_12871_),
    .Y(_12872_));
 sky130_fd_sc_hd__o22ai_1 _18743_ (.A1(net3524),
    .A2(_12870_),
    .B1(_12872_),
    .B2(_12394_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand3_2 _18744_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(\cs_registers_i.pc_id_i[24] ),
    .C(_12863_),
    .Y(_12873_));
 sky130_fd_sc_hd__xnor2_1 _18745_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(_12873_),
    .Y(_12874_));
 sky130_fd_sc_hd__a222oi_1 _18746_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net3609),
    .B1(_12874_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net379),
    .Y(_12875_));
 sky130_fd_sc_hd__nor2_1 _18747_ (.A(_11457_),
    .B(_12757_),
    .Y(_12876_));
 sky130_fd_sc_hd__a21oi_1 _18748_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_12757_),
    .B1(_12876_),
    .Y(_12877_));
 sky130_fd_sc_hd__o22ai_1 _18749_ (.A1(net3524),
    .A2(_12875_),
    .B1(_12877_),
    .B2(net3532),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_1 _18750_ (.A(\cs_registers_i.pc_id_i[25] ),
    .Y(_12878_));
 sky130_fd_sc_hd__nor2_2 _18751_ (.A(_12878_),
    .B(_12873_),
    .Y(_12879_));
 sky130_fd_sc_hd__xor2_1 _18752_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(_12879_),
    .X(_12880_));
 sky130_fd_sc_hd__a222oi_1 _18753_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net3609),
    .B1(_12880_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3842),
    .Y(_12881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_656 ();
 sky130_fd_sc_hd__nor2_1 _18755_ (.A(_11476_),
    .B(_12757_),
    .Y(_12883_));
 sky130_fd_sc_hd__a21oi_1 _18756_ (.A1(\cs_registers_i.mtval_q[26] ),
    .A2(_12757_),
    .B1(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__o22ai_1 _18757_ (.A1(net3524),
    .A2(_12881_),
    .B1(_12884_),
    .B2(net3532),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _18758_ (.A(net3826),
    .B(_12879_),
    .Y(_12885_));
 sky130_fd_sc_hd__xnor2_1 _18759_ (.A(net3825),
    .B(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__a222oi_1 _18760_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net3609),
    .B1(_12886_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3841),
    .Y(_12887_));
 sky130_fd_sc_hd__nor2_1 _18761_ (.A(_11490_),
    .B(_12757_),
    .Y(_12888_));
 sky130_fd_sc_hd__a21oi_1 _18762_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(_12757_),
    .B1(_12888_),
    .Y(_12889_));
 sky130_fd_sc_hd__o22ai_1 _18763_ (.A1(net3524),
    .A2(_12887_),
    .B1(_12889_),
    .B2(net3532),
    .Y(_00406_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_655 ();
 sky130_fd_sc_hd__nand3_2 _18765_ (.A(net3826),
    .B(\cs_registers_i.pc_id_i[27] ),
    .C(_12879_),
    .Y(_12891_));
 sky130_fd_sc_hd__xnor2_1 _18766_ (.A(net3824),
    .B(_12891_),
    .Y(_12892_));
 sky130_fd_sc_hd__a222oi_1 _18767_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net3609),
    .B1(_12892_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net368),
    .Y(_12893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_654 ();
 sky130_fd_sc_hd__nor2_1 _18769_ (.A(_11506_),
    .B(_12757_),
    .Y(_12895_));
 sky130_fd_sc_hd__a21oi_1 _18770_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(_12757_),
    .B1(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_653 ();
 sky130_fd_sc_hd__o22ai_1 _18772_ (.A1(net3524),
    .A2(_12893_),
    .B1(_12896_),
    .B2(_12394_),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_1 _18773_ (.A(net3824),
    .Y(_12898_));
 sky130_fd_sc_hd__nor2_2 _18774_ (.A(_12898_),
    .B(_12891_),
    .Y(_12899_));
 sky130_fd_sc_hd__xor2_1 _18775_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_12899_),
    .X(_12900_));
 sky130_fd_sc_hd__a222oi_1 _18776_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net3609),
    .B1(_12900_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3839),
    .Y(_12901_));
 sky130_fd_sc_hd__nor2_1 _18777_ (.A(_11530_),
    .B(_12757_),
    .Y(_12902_));
 sky130_fd_sc_hd__a21oi_1 _18778_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_12757_),
    .B1(_12902_),
    .Y(_12903_));
 sky130_fd_sc_hd__o22ai_1 _18779_ (.A1(net3524),
    .A2(_12901_),
    .B1(_12903_),
    .B2(_12394_),
    .Y(_00408_));
 sky130_fd_sc_hd__xnor2_1 _18780_ (.A(_08414_),
    .B(_12765_),
    .Y(_12904_));
 sky130_fd_sc_hd__mux2i_1 _18781_ (.A0(net338),
    .A1(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .S(net3947),
    .Y(_12905_));
 sky130_fd_sc_hd__o22ai_1 _18782_ (.A1(_10646_),
    .A2(_12904_),
    .B1(_12905_),
    .B2(_12748_),
    .Y(_12906_));
 sky130_fd_sc_hd__a21oi_2 _18783_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(net3609),
    .B1(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__nor2_1 _18784_ (.A(_11082_),
    .B(_12757_),
    .Y(_12908_));
 sky130_fd_sc_hd__a21oi_1 _18785_ (.A1(\cs_registers_i.mtval_q[2] ),
    .A2(_12757_),
    .B1(_12908_),
    .Y(_12909_));
 sky130_fd_sc_hd__o22ai_1 _18786_ (.A1(net3524),
    .A2(_12907_),
    .B1(_12909_),
    .B2(_12394_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _18787_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_12899_),
    .Y(_12910_));
 sky130_fd_sc_hd__xnor2_1 _18788_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__a222oi_1 _18789_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net3609),
    .B1(_12911_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net354),
    .Y(_12912_));
 sky130_fd_sc_hd__nor2_1 _18790_ (.A(_11550_),
    .B(_12757_),
    .Y(_12913_));
 sky130_fd_sc_hd__a21oi_1 _18791_ (.A1(\cs_registers_i.mtval_q[30] ),
    .A2(_12757_),
    .B1(_12913_),
    .Y(_12914_));
 sky130_fd_sc_hd__o22ai_1 _18792_ (.A1(net3524),
    .A2(_12912_),
    .B1(_12914_),
    .B2(net3532),
    .Y(_00410_));
 sky130_fd_sc_hd__nand3_1 _18793_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(\cs_registers_i.pc_id_i[30] ),
    .C(_12899_),
    .Y(_12915_));
 sky130_fd_sc_hd__xnor2_1 _18794_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(_12915_),
    .Y(_12916_));
 sky130_fd_sc_hd__a222oi_1 _18795_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net3609),
    .B1(_12916_),
    .B2(_12416_),
    .C1(_12813_),
    .C2(net3836),
    .Y(_12917_));
 sky130_fd_sc_hd__nor2_1 _18796_ (.A(_11565_),
    .B(_12757_),
    .Y(_12918_));
 sky130_fd_sc_hd__a21oi_1 _18797_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(_12757_),
    .B1(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__o22ai_1 _18798_ (.A1(net3524),
    .A2(_12917_),
    .B1(_12919_),
    .B2(_12394_),
    .Y(_00411_));
 sky130_fd_sc_hd__a31oi_1 _18799_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .B1(\cs_registers_i.pc_id_i[3] ),
    .Y(_12920_));
 sky130_fd_sc_hd__mux2i_1 _18800_ (.A0(net3835),
    .A1(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .S(net3947),
    .Y(_12921_));
 sky130_fd_sc_hd__o32ai_2 _18801_ (.A1(_10646_),
    .A2(_12766_),
    .A3(_12920_),
    .B1(_12921_),
    .B2(_12748_),
    .Y(_12922_));
 sky130_fd_sc_hd__a21oi_4 _18802_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(net3609),
    .B1(_12922_),
    .Y(_12923_));
 sky130_fd_sc_hd__nor2_1 _18803_ (.A(_11612_),
    .B(_12757_),
    .Y(_12924_));
 sky130_fd_sc_hd__a21oi_1 _18804_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(_12757_),
    .B1(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__o22ai_1 _18805_ (.A1(net3524),
    .A2(_12923_),
    .B1(_12925_),
    .B2(net3532),
    .Y(_00412_));
 sky130_fd_sc_hd__mux2i_1 _18806_ (.A0(net325),
    .A1(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .S(net3947),
    .Y(_12926_));
 sky130_fd_sc_hd__xnor2_1 _18807_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(_12766_),
    .Y(_12927_));
 sky130_fd_sc_hd__o22ai_1 _18808_ (.A1(_12748_),
    .A2(_12926_),
    .B1(_12927_),
    .B2(_10646_),
    .Y(_12928_));
 sky130_fd_sc_hd__a21oi_1 _18809_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(net3609),
    .B1(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__nor2_1 _18810_ (.A(_11780_),
    .B(_12757_),
    .Y(_12930_));
 sky130_fd_sc_hd__a21oi_1 _18811_ (.A1(\cs_registers_i.mtval_q[4] ),
    .A2(_12757_),
    .B1(_12930_),
    .Y(_12931_));
 sky130_fd_sc_hd__o22ai_1 _18812_ (.A1(net3524),
    .A2(_12929_),
    .B1(_12931_),
    .B2(_12394_),
    .Y(_00413_));
 sky130_fd_sc_hd__a21oi_1 _18813_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_12766_),
    .B1(\cs_registers_i.pc_id_i[5] ),
    .Y(_12932_));
 sky130_fd_sc_hd__mux2i_1 _18814_ (.A0(net3831),
    .A1(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .S(net3947),
    .Y(_12933_));
 sky130_fd_sc_hd__o32ai_2 _18815_ (.A1(_10646_),
    .A2(_12767_),
    .A3(_12932_),
    .B1(_12933_),
    .B2(_12748_),
    .Y(_12934_));
 sky130_fd_sc_hd__a21oi_1 _18816_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(net3609),
    .B1(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__nor2_1 _18817_ (.A(_11647_),
    .B(_12757_),
    .Y(_12936_));
 sky130_fd_sc_hd__a21oi_1 _18818_ (.A1(\cs_registers_i.mtval_q[5] ),
    .A2(_12757_),
    .B1(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__o22ai_1 _18819_ (.A1(net3524),
    .A2(_12935_),
    .B1(_12937_),
    .B2(_12394_),
    .Y(_00414_));
 sky130_fd_sc_hd__mux2i_1 _18820_ (.A0(\id_stage_i.controller_i.instr_i[6] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .S(net3947),
    .Y(_12938_));
 sky130_fd_sc_hd__xnor2_1 _18821_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(_12767_),
    .Y(_12939_));
 sky130_fd_sc_hd__o22ai_1 _18822_ (.A1(_12748_),
    .A2(_12938_),
    .B1(_12939_),
    .B2(_10646_),
    .Y(_12940_));
 sky130_fd_sc_hd__a21oi_1 _18823_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net3609),
    .B1(_12940_),
    .Y(_12941_));
 sky130_fd_sc_hd__nor2_1 _18824_ (.A(_11664_),
    .B(_12757_),
    .Y(_12942_));
 sky130_fd_sc_hd__a21oi_1 _18825_ (.A1(\cs_registers_i.mtval_q[6] ),
    .A2(_12757_),
    .B1(_12942_),
    .Y(_12943_));
 sky130_fd_sc_hd__o22ai_1 _18826_ (.A1(net3524),
    .A2(_12941_),
    .B1(_12943_),
    .B2(_12394_),
    .Y(_00415_));
 sky130_fd_sc_hd__a21oi_1 _18827_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_12767_),
    .B1(\cs_registers_i.pc_id_i[7] ),
    .Y(_12944_));
 sky130_fd_sc_hd__mux2i_2 _18828_ (.A0(net3829),
    .A1(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .S(net3947),
    .Y(_12945_));
 sky130_fd_sc_hd__o32ai_1 _18829_ (.A1(_10646_),
    .A2(_12768_),
    .A3(_12944_),
    .B1(_12945_),
    .B2(_12748_),
    .Y(_12946_));
 sky130_fd_sc_hd__a21oi_1 _18830_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net3609),
    .B1(_12946_),
    .Y(_12947_));
 sky130_fd_sc_hd__nor2_1 _18831_ (.A(_11685_),
    .B(_12757_),
    .Y(_12948_));
 sky130_fd_sc_hd__a21oi_1 _18832_ (.A1(\cs_registers_i.mtval_q[7] ),
    .A2(_12757_),
    .B1(_12948_),
    .Y(_12949_));
 sky130_fd_sc_hd__o22ai_1 _18833_ (.A1(net3524),
    .A2(_12947_),
    .B1(_12949_),
    .B2(_12394_),
    .Y(_00416_));
 sky130_fd_sc_hd__mux2i_2 _18834_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .S(net3947),
    .Y(_12950_));
 sky130_fd_sc_hd__xnor2_1 _18835_ (.A(net3823),
    .B(_12768_),
    .Y(_12951_));
 sky130_fd_sc_hd__o22ai_1 _18836_ (.A1(_12748_),
    .A2(_12950_),
    .B1(_12951_),
    .B2(_10646_),
    .Y(_12952_));
 sky130_fd_sc_hd__a21oi_2 _18837_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(net3609),
    .B1(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__nor2_1 _18838_ (.A(_11707_),
    .B(_12757_),
    .Y(_12954_));
 sky130_fd_sc_hd__a21oi_1 _18839_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(_12757_),
    .B1(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__o22ai_1 _18840_ (.A1(net3524),
    .A2(_12953_),
    .B1(_12955_),
    .B2(_12394_),
    .Y(_00417_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_652 ();
 sky130_fd_sc_hd__mux2_8 _18842_ (.A0(net3827),
    .A1(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .S(net3947),
    .X(_12957_));
 sky130_fd_sc_hd__nand2_1 _18843_ (.A(net3823),
    .B(_12768_),
    .Y(_12958_));
 sky130_fd_sc_hd__xnor2_1 _18844_ (.A(\cs_registers_i.pc_id_i[9] ),
    .B(_12958_),
    .Y(_12959_));
 sky130_fd_sc_hd__a222oi_1 _18845_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(net3609),
    .B1(_12452_),
    .B2(_12957_),
    .C1(_12959_),
    .C2(_12416_),
    .Y(_12960_));
 sky130_fd_sc_hd__nor2_1 _18846_ (.A(_11726_),
    .B(_12757_),
    .Y(_12961_));
 sky130_fd_sc_hd__a21oi_1 _18847_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(_12757_),
    .B1(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__o22ai_1 _18848_ (.A1(net3524),
    .A2(_12960_),
    .B1(_12962_),
    .B2(_12394_),
    .Y(_00418_));
 sky130_fd_sc_hd__or3_4 _18849_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .X(_12963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_650 ();
 sky130_fd_sc_hd__nand2_8 _18852_ (.A(net3550),
    .B(net3501),
    .Y(_12966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_647 ();
 sky130_fd_sc_hd__nor2_1 _18856_ (.A(_11145_),
    .B(_12966_),
    .Y(_12970_));
 sky130_fd_sc_hd__a21oi_1 _18857_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(_12966_),
    .B1(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_646 ();
 sky130_fd_sc_hd__nor2_1 _18859_ (.A(net1),
    .B(_12963_),
    .Y(_12973_));
 sky130_fd_sc_hd__a21oi_1 _18860_ (.A1(_12963_),
    .A2(_12971_),
    .B1(_12973_),
    .Y(_00419_));
 sky130_fd_sc_hd__nor2_1 _18861_ (.A(_11177_),
    .B(_12966_),
    .Y(_12974_));
 sky130_fd_sc_hd__a21oi_1 _18862_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_12966_),
    .B1(_12974_),
    .Y(_12975_));
 sky130_fd_sc_hd__nor2_1 _18863_ (.A(net2),
    .B(_12963_),
    .Y(_12976_));
 sky130_fd_sc_hd__a21oi_1 _18864_ (.A1(_12963_),
    .A2(_12975_),
    .B1(_12976_),
    .Y(_00420_));
 sky130_fd_sc_hd__nor2_1 _18865_ (.A(_11197_),
    .B(_12966_),
    .Y(_12977_));
 sky130_fd_sc_hd__a21oi_1 _18866_ (.A1(\cs_registers_i.csr_mtvec_o[12] ),
    .A2(_12966_),
    .B1(_12977_),
    .Y(_12978_));
 sky130_fd_sc_hd__nor2_1 _18867_ (.A(net3),
    .B(_12963_),
    .Y(_12979_));
 sky130_fd_sc_hd__a21oi_1 _18868_ (.A1(_12963_),
    .A2(_12978_),
    .B1(_12979_),
    .Y(_00421_));
 sky130_fd_sc_hd__nor2_1 _18869_ (.A(_11214_),
    .B(_12966_),
    .Y(_12980_));
 sky130_fd_sc_hd__a21oi_1 _18870_ (.A1(\cs_registers_i.csr_mtvec_o[13] ),
    .A2(_12966_),
    .B1(_12980_),
    .Y(_12981_));
 sky130_fd_sc_hd__nor2_1 _18871_ (.A(net4),
    .B(_12963_),
    .Y(_12982_));
 sky130_fd_sc_hd__a21oi_1 _18872_ (.A1(_12963_),
    .A2(_12981_),
    .B1(_12982_),
    .Y(_00422_));
 sky130_fd_sc_hd__nor2_1 _18873_ (.A(_11235_),
    .B(_12966_),
    .Y(_12983_));
 sky130_fd_sc_hd__a21oi_1 _18874_ (.A1(\cs_registers_i.csr_mtvec_o[14] ),
    .A2(_12966_),
    .B1(_12983_),
    .Y(_12984_));
 sky130_fd_sc_hd__nor2_1 _18875_ (.A(net5),
    .B(_12963_),
    .Y(_12985_));
 sky130_fd_sc_hd__a21oi_1 _18876_ (.A1(_12963_),
    .A2(_12984_),
    .B1(_12985_),
    .Y(_00423_));
 sky130_fd_sc_hd__nor2_1 _18877_ (.A(_11255_),
    .B(_12966_),
    .Y(_12986_));
 sky130_fd_sc_hd__a21oi_1 _18878_ (.A1(\cs_registers_i.csr_mtvec_o[15] ),
    .A2(_12966_),
    .B1(_12986_),
    .Y(_12987_));
 sky130_fd_sc_hd__nor2_1 _18879_ (.A(net6),
    .B(_12963_),
    .Y(_12988_));
 sky130_fd_sc_hd__a21oi_1 _18880_ (.A1(_12963_),
    .A2(_12987_),
    .B1(_12988_),
    .Y(_00424_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_645 ();
 sky130_fd_sc_hd__nor2_1 _18882_ (.A(_11270_),
    .B(_12966_),
    .Y(_12990_));
 sky130_fd_sc_hd__a21oi_1 _18883_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_12966_),
    .B1(_12990_),
    .Y(_12991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_644 ();
 sky130_fd_sc_hd__nor2_1 _18885_ (.A(net7),
    .B(_12963_),
    .Y(_12993_));
 sky130_fd_sc_hd__a21oi_1 _18886_ (.A1(_12963_),
    .A2(_12991_),
    .B1(_12993_),
    .Y(_00425_));
 sky130_fd_sc_hd__nor2_1 _18887_ (.A(_11294_),
    .B(_12966_),
    .Y(_12994_));
 sky130_fd_sc_hd__a21oi_1 _18888_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(_12966_),
    .B1(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__nor2_1 _18889_ (.A(net8),
    .B(_12963_),
    .Y(_12996_));
 sky130_fd_sc_hd__a21oi_1 _18890_ (.A1(_12963_),
    .A2(_12995_),
    .B1(_12996_),
    .Y(_00426_));
 sky130_fd_sc_hd__nor2_1 _18891_ (.A(_11319_),
    .B(_12966_),
    .Y(_12997_));
 sky130_fd_sc_hd__a21oi_1 _18892_ (.A1(\cs_registers_i.csr_mtvec_o[18] ),
    .A2(_12966_),
    .B1(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__nor2_1 _18893_ (.A(net9),
    .B(_12963_),
    .Y(_12999_));
 sky130_fd_sc_hd__a21oi_1 _18894_ (.A1(_12963_),
    .A2(_12998_),
    .B1(_12999_),
    .Y(_00427_));
 sky130_fd_sc_hd__nor2_1 _18895_ (.A(_11333_),
    .B(_12966_),
    .Y(_13000_));
 sky130_fd_sc_hd__a21oi_1 _18896_ (.A1(\cs_registers_i.csr_mtvec_o[19] ),
    .A2(_12966_),
    .B1(_13000_),
    .Y(_13001_));
 sky130_fd_sc_hd__nor2_1 _18897_ (.A(net10),
    .B(_12963_),
    .Y(_13002_));
 sky130_fd_sc_hd__a21oi_1 _18898_ (.A1(_12963_),
    .A2(_13001_),
    .B1(_13002_),
    .Y(_00428_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_642 ();
 sky130_fd_sc_hd__nor2_1 _18901_ (.A(_11369_),
    .B(_12966_),
    .Y(_13005_));
 sky130_fd_sc_hd__a21oi_1 _18902_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_12966_),
    .B1(_13005_),
    .Y(_13006_));
 sky130_fd_sc_hd__nor2_1 _18903_ (.A(net11),
    .B(_12963_),
    .Y(_13007_));
 sky130_fd_sc_hd__a21oi_1 _18904_ (.A1(_12963_),
    .A2(_13006_),
    .B1(_13007_),
    .Y(_00429_));
 sky130_fd_sc_hd__nor2_1 _18905_ (.A(_11390_),
    .B(_12966_),
    .Y(_13008_));
 sky130_fd_sc_hd__a21oi_1 _18906_ (.A1(\cs_registers_i.csr_mtvec_o[21] ),
    .A2(_12966_),
    .B1(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__nor2_1 _18907_ (.A(net12),
    .B(_12963_),
    .Y(_13010_));
 sky130_fd_sc_hd__a21oi_1 _18908_ (.A1(_12963_),
    .A2(_13009_),
    .B1(_13010_),
    .Y(_00430_));
 sky130_fd_sc_hd__nor2_1 _18909_ (.A(_11406_),
    .B(_12966_),
    .Y(_13011_));
 sky130_fd_sc_hd__a21oi_1 _18910_ (.A1(\cs_registers_i.csr_mtvec_o[22] ),
    .A2(_12966_),
    .B1(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__nor2_1 _18911_ (.A(net13),
    .B(_12963_),
    .Y(_13013_));
 sky130_fd_sc_hd__a21oi_1 _18912_ (.A1(_12963_),
    .A2(_13012_),
    .B1(_13013_),
    .Y(_00431_));
 sky130_fd_sc_hd__nor2_1 _18913_ (.A(_11426_),
    .B(_12966_),
    .Y(_13014_));
 sky130_fd_sc_hd__a21oi_1 _18914_ (.A1(\cs_registers_i.csr_mtvec_o[23] ),
    .A2(_12966_),
    .B1(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__nor2_1 _18915_ (.A(net14),
    .B(_12963_),
    .Y(_13016_));
 sky130_fd_sc_hd__a21oi_1 _18916_ (.A1(_12963_),
    .A2(_13015_),
    .B1(_13016_),
    .Y(_00432_));
 sky130_fd_sc_hd__nor2_1 _18917_ (.A(_11441_),
    .B(_12966_),
    .Y(_13017_));
 sky130_fd_sc_hd__a21oi_1 _18918_ (.A1(\cs_registers_i.csr_mtvec_o[24] ),
    .A2(_12966_),
    .B1(_13017_),
    .Y(_13018_));
 sky130_fd_sc_hd__nor2_1 _18919_ (.A(net15),
    .B(_12963_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21oi_1 _18920_ (.A1(_12963_),
    .A2(_13018_),
    .B1(_13019_),
    .Y(_00433_));
 sky130_fd_sc_hd__nor2_1 _18921_ (.A(_11457_),
    .B(_12966_),
    .Y(_13020_));
 sky130_fd_sc_hd__a21oi_1 _18922_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_12966_),
    .B1(_13020_),
    .Y(_13021_));
 sky130_fd_sc_hd__nor2_1 _18923_ (.A(net16),
    .B(_12963_),
    .Y(_13022_));
 sky130_fd_sc_hd__a21oi_1 _18924_ (.A1(_12963_),
    .A2(_13021_),
    .B1(_13022_),
    .Y(_00434_));
 sky130_fd_sc_hd__nor2_1 _18925_ (.A(_11476_),
    .B(_12966_),
    .Y(_13023_));
 sky130_fd_sc_hd__a21oi_1 _18926_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(_12966_),
    .B1(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__nor2_1 _18927_ (.A(net17),
    .B(_12963_),
    .Y(_13025_));
 sky130_fd_sc_hd__a21oi_1 _18928_ (.A1(_12963_),
    .A2(_13024_),
    .B1(_13025_),
    .Y(_00435_));
 sky130_fd_sc_hd__nor2_1 _18929_ (.A(_11490_),
    .B(_12966_),
    .Y(_13026_));
 sky130_fd_sc_hd__a21oi_1 _18930_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_12966_),
    .B1(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__nor2_1 _18931_ (.A(net18),
    .B(_12963_),
    .Y(_13028_));
 sky130_fd_sc_hd__a21oi_1 _18932_ (.A1(_12963_),
    .A2(_13027_),
    .B1(_13028_),
    .Y(_00436_));
 sky130_fd_sc_hd__nor2_1 _18933_ (.A(_11506_),
    .B(_12966_),
    .Y(_13029_));
 sky130_fd_sc_hd__a21oi_1 _18934_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_12966_),
    .B1(_13029_),
    .Y(_13030_));
 sky130_fd_sc_hd__nor2_1 _18935_ (.A(net19),
    .B(_12963_),
    .Y(_13031_));
 sky130_fd_sc_hd__a21oi_1 _18936_ (.A1(_12963_),
    .A2(_13030_),
    .B1(_13031_),
    .Y(_00437_));
 sky130_fd_sc_hd__nor2_1 _18937_ (.A(_11530_),
    .B(_12966_),
    .Y(_13032_));
 sky130_fd_sc_hd__a21oi_1 _18938_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(_12966_),
    .B1(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__nor2_1 _18939_ (.A(net20),
    .B(_12963_),
    .Y(_13034_));
 sky130_fd_sc_hd__a21oi_1 _18940_ (.A1(_12963_),
    .A2(_13033_),
    .B1(_13034_),
    .Y(_00438_));
 sky130_fd_sc_hd__nor2_1 _18941_ (.A(_11550_),
    .B(_12966_),
    .Y(_13035_));
 sky130_fd_sc_hd__a21oi_1 _18942_ (.A1(\cs_registers_i.csr_mtvec_o[30] ),
    .A2(_12966_),
    .B1(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__nor2_1 _18943_ (.A(net21),
    .B(_12963_),
    .Y(_13037_));
 sky130_fd_sc_hd__a21oi_1 _18944_ (.A1(_12963_),
    .A2(_13036_),
    .B1(_13037_),
    .Y(_00439_));
 sky130_fd_sc_hd__nor2_1 _18945_ (.A(_11565_),
    .B(_12966_),
    .Y(_13038_));
 sky130_fd_sc_hd__a21oi_1 _18946_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_12966_),
    .B1(_13038_),
    .Y(_13039_));
 sky130_fd_sc_hd__nor2_1 _18947_ (.A(net22),
    .B(_12963_),
    .Y(_13040_));
 sky130_fd_sc_hd__a21oi_1 _18948_ (.A1(_12963_),
    .A2(_13039_),
    .B1(_13040_),
    .Y(_00440_));
 sky130_fd_sc_hd__nor2_1 _18949_ (.A(_11707_),
    .B(_12966_),
    .Y(_13041_));
 sky130_fd_sc_hd__a21oi_1 _18950_ (.A1(\cs_registers_i.csr_mtvec_o[8] ),
    .A2(_12966_),
    .B1(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__nor2_1 _18951_ (.A(net23),
    .B(_12963_),
    .Y(_13043_));
 sky130_fd_sc_hd__a21oi_1 _18952_ (.A1(_12963_),
    .A2(_13042_),
    .B1(_13043_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2_1 _18953_ (.A(_11726_),
    .B(_12966_),
    .Y(_13044_));
 sky130_fd_sc_hd__a21oi_1 _18954_ (.A1(\cs_registers_i.csr_mtvec_o[9] ),
    .A2(_12966_),
    .B1(_13044_),
    .Y(_13045_));
 sky130_fd_sc_hd__nor2_1 _18955_ (.A(net24),
    .B(_12963_),
    .Y(_13046_));
 sky130_fd_sc_hd__a21oi_1 _18956_ (.A1(_12963_),
    .A2(_13045_),
    .B1(_13046_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_8 _18957_ (.A(net3936),
    .B(_07857_),
    .Y(_13047_));
 sky130_fd_sc_hd__nor2_4 _18958_ (.A(net3940),
    .B(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_640 ();
 sky130_fd_sc_hd__nand3_1 _18961_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .B(_10980_),
    .C(_13048_),
    .Y(_13051_));
 sky130_fd_sc_hd__mux2_1 _18962_ (.A0(_10736_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .S(_13051_),
    .X(_00443_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_638 ();
 sky130_fd_sc_hd__nor3_2 _18965_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .Y(_13054_));
 sky130_fd_sc_hd__and2_4 _18966_ (.A(_10980_),
    .B(_13054_),
    .X(_13055_));
 sky130_fd_sc_hd__nor2_1 _18967_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_10980_),
    .Y(_13056_));
 sky130_fd_sc_hd__a21oi_1 _18968_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A2(_13055_),
    .B1(_13056_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_4 _18969_ (.A(_10672_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_13057_));
 sky130_fd_sc_hd__nand2_1 _18970_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_13054_),
    .Y(_13058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_637 ();
 sky130_fd_sc_hd__a21oi_1 _18972_ (.A1(_10980_),
    .A2(_13058_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_13060_));
 sky130_fd_sc_hd__a21oi_1 _18973_ (.A1(_13055_),
    .A2(_13057_),
    .B1(_13060_),
    .Y(_00445_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_636 ();
 sky130_fd_sc_hd__nor2_1 _18975_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_13062_));
 sky130_fd_sc_hd__and2_4 _18976_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13062_),
    .X(_13063_));
 sky130_fd_sc_hd__o21ai_0 _18977_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B1(_13054_),
    .Y(_13064_));
 sky130_fd_sc_hd__a21oi_1 _18978_ (.A1(_10980_),
    .A2(_13064_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13065_));
 sky130_fd_sc_hd__a21oi_1 _18979_ (.A1(_13055_),
    .A2(_13063_),
    .B1(_13065_),
    .Y(_00446_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_635 ();
 sky130_fd_sc_hd__nor3_2 _18981_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13067_));
 sky130_fd_sc_hd__or3_4 _18982_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .X(_13068_));
 sky130_fd_sc_hd__nand2_1 _18983_ (.A(_13054_),
    .B(_13068_),
    .Y(_13069_));
 sky130_fd_sc_hd__a21oi_1 _18984_ (.A1(_10980_),
    .A2(_13069_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .Y(_13070_));
 sky130_fd_sc_hd__a31oi_1 _18985_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_13055_),
    .A3(_13067_),
    .B1(_13070_),
    .Y(_00447_));
 sky130_fd_sc_hd__nor2_4 _18986_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_13068_),
    .Y(_13071_));
 sky130_fd_sc_hd__o21ai_0 _18987_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_13068_),
    .B1(_13054_),
    .Y(_13072_));
 sky130_fd_sc_hd__a21oi_1 _18988_ (.A1(_10980_),
    .A2(_13072_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .Y(_13073_));
 sky130_fd_sc_hd__a31oi_1 _18989_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_13055_),
    .A3(_13071_),
    .B1(_13073_),
    .Y(_00448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_634 ();
 sky130_fd_sc_hd__o21ai_2 _18991_ (.A1(net3939),
    .A2(net3936),
    .B1(net3944),
    .Y(_13075_));
 sky130_fd_sc_hd__nand2_8 _18992_ (.A(_08075_),
    .B(_13075_),
    .Y(_13076_));
 sky130_fd_sc_hd__nor2_2 _18993_ (.A(net321),
    .B(_13076_),
    .Y(_13077_));
 sky130_fd_sc_hd__and4_4 _18994_ (.A(_10402_),
    .B(_10409_),
    .C(_10414_),
    .D(_13077_),
    .X(_13078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_633 ();
 sky130_fd_sc_hd__mux2_1 _18996_ (.A0(net3711),
    .A1(net3575),
    .S(net3672),
    .X(_13080_));
 sky130_fd_sc_hd__nand2_8 _18997_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(_10980_),
    .Y(_13081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_632 ();
 sky130_fd_sc_hd__nand2_1 _18999_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .B(_13081_),
    .Y(_13083_));
 sky130_fd_sc_hd__o21ai_0 _19000_ (.A1(_10984_),
    .A2(_13080_),
    .B1(_13083_),
    .Y(_00449_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_630 ();
 sky130_fd_sc_hd__nor2_1 _19003_ (.A(net400),
    .B(net3672),
    .Y(_13086_));
 sky130_fd_sc_hd__a21oi_1 _19004_ (.A1(net151),
    .A2(net3672),
    .B1(_13086_),
    .Y(_13087_));
 sky130_fd_sc_hd__nand2_1 _19005_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .B(_13081_),
    .Y(_13088_));
 sky130_fd_sc_hd__o21ai_0 _19006_ (.A1(_10984_),
    .A2(_13087_),
    .B1(_13088_),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_1 _19007_ (.A(net3703),
    .B(net3672),
    .Y(_13089_));
 sky130_fd_sc_hd__a21oi_1 _19008_ (.A1(net152),
    .A2(net3672),
    .B1(_13089_),
    .Y(_13090_));
 sky130_fd_sc_hd__nand2_1 _19009_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .B(_13081_),
    .Y(_13091_));
 sky130_fd_sc_hd__o21ai_0 _19010_ (.A1(_10984_),
    .A2(_13090_),
    .B1(_13091_),
    .Y(_00451_));
 sky130_fd_sc_hd__nor2_1 _19011_ (.A(net401),
    .B(net3672),
    .Y(_13092_));
 sky130_fd_sc_hd__a21oi_1 _19012_ (.A1(net3514),
    .A2(net3672),
    .B1(_13092_),
    .Y(_13093_));
 sky130_fd_sc_hd__nand2_1 _19013_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .B(_13081_),
    .Y(_13094_));
 sky130_fd_sc_hd__o21ai_0 _19014_ (.A1(_10984_),
    .A2(_13093_),
    .B1(_13094_),
    .Y(_00452_));
 sky130_fd_sc_hd__nor2_1 _19015_ (.A(net3699),
    .B(net3672),
    .Y(_13095_));
 sky130_fd_sc_hd__a21oi_1 _19016_ (.A1(net154),
    .A2(net3672),
    .B1(_13095_),
    .Y(_13096_));
 sky130_fd_sc_hd__nand2_1 _19017_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .B(_13081_),
    .Y(_13097_));
 sky130_fd_sc_hd__o21ai_0 _19018_ (.A1(_10984_),
    .A2(_13096_),
    .B1(_13097_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand4_4 _19019_ (.A(_10402_),
    .B(_10409_),
    .C(_10414_),
    .D(_13077_),
    .Y(_13098_));
 sky130_fd_sc_hd__nand2_1 _19020_ (.A(net3695),
    .B(_13098_),
    .Y(_13099_));
 sky130_fd_sc_hd__o21ai_1 _19021_ (.A1(net3513),
    .A2(_13098_),
    .B1(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_1 _19022_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .B(_13081_),
    .Y(_13101_));
 sky130_fd_sc_hd__o21ai_0 _19023_ (.A1(_10984_),
    .A2(_13100_),
    .B1(_13101_),
    .Y(_00454_));
 sky130_fd_sc_hd__nor2_1 _19024_ (.A(net3697),
    .B(net3672),
    .Y(_13102_));
 sky130_fd_sc_hd__a21oi_2 _19025_ (.A1(net3507),
    .A2(net3672),
    .B1(_13102_),
    .Y(_13103_));
 sky130_fd_sc_hd__nand2_1 _19026_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .B(_13081_),
    .Y(_13104_));
 sky130_fd_sc_hd__o21ai_0 _19027_ (.A1(_10984_),
    .A2(_13103_),
    .B1(_13104_),
    .Y(_00455_));
 sky130_fd_sc_hd__nor2_1 _19028_ (.A(net3693),
    .B(_13078_),
    .Y(_13105_));
 sky130_fd_sc_hd__a21oi_1 _19029_ (.A1(net3506),
    .A2(_13078_),
    .B1(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__nand2_1 _19030_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .B(_13081_),
    .Y(_13107_));
 sky130_fd_sc_hd__o21ai_0 _19031_ (.A1(_10984_),
    .A2(_13106_),
    .B1(_13107_),
    .Y(_00456_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_629 ();
 sky130_fd_sc_hd__mux2i_1 _19033_ (.A0(net332),
    .A1(net420),
    .S(_13078_),
    .Y(_13109_));
 sky130_fd_sc_hd__nand2_1 _19034_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .B(_13081_),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ai_0 _19035_ (.A1(_10984_),
    .A2(_13109_),
    .B1(_13110_),
    .Y(_00457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_628 ();
 sky130_fd_sc_hd__nor2_1 _19037_ (.A(_09652_),
    .B(_13078_),
    .Y(_13112_));
 sky130_fd_sc_hd__a21oi_1 _19038_ (.A1(net159),
    .A2(_13078_),
    .B1(_13112_),
    .Y(_13113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_627 ();
 sky130_fd_sc_hd__nand2_1 _19040_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .B(_13081_),
    .Y(_13115_));
 sky130_fd_sc_hd__o21ai_0 _19041_ (.A1(_10984_),
    .A2(_13113_),
    .B1(_13115_),
    .Y(_00458_));
 sky130_fd_sc_hd__mux2i_1 _19042_ (.A0(net422),
    .A1(net160),
    .S(_13078_),
    .Y(_13116_));
 sky130_fd_sc_hd__nand2_1 _19043_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .B(_13081_),
    .Y(_13117_));
 sky130_fd_sc_hd__o21ai_0 _19044_ (.A1(_10984_),
    .A2(_13116_),
    .B1(_13117_),
    .Y(_00459_));
 sky130_fd_sc_hd__xor2_4 _19045_ (.A(net3583),
    .B(net3574),
    .X(_13118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_626 ();
 sky130_fd_sc_hd__nor2_1 _19047_ (.A(_13098_),
    .B(_13118_),
    .Y(_13120_));
 sky130_fd_sc_hd__a21oi_2 _19048_ (.A1(net3714),
    .A2(_13098_),
    .B1(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__nand2_1 _19049_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .B(_13081_),
    .Y(_13122_));
 sky130_fd_sc_hd__o21ai_0 _19050_ (.A1(_10984_),
    .A2(_13121_),
    .B1(_13122_),
    .Y(_00460_));
 sky130_fd_sc_hd__nor2_1 _19051_ (.A(net3689),
    .B(_13078_),
    .Y(_13123_));
 sky130_fd_sc_hd__a21oi_1 _19052_ (.A1(net452),
    .A2(_13078_),
    .B1(_13123_),
    .Y(_13124_));
 sky130_fd_sc_hd__nand2_1 _19053_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .B(_13081_),
    .Y(_13125_));
 sky130_fd_sc_hd__o21ai_0 _19054_ (.A1(_10984_),
    .A2(_13124_),
    .B1(_13125_),
    .Y(_00461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_625 ();
 sky130_fd_sc_hd__nor2_1 _19056_ (.A(net3690),
    .B(_13078_),
    .Y(_13127_));
 sky130_fd_sc_hd__a21oi_1 _19057_ (.A1(net162),
    .A2(_13078_),
    .B1(_13127_),
    .Y(_13128_));
 sky130_fd_sc_hd__nand2_1 _19058_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .B(_13081_),
    .Y(_13129_));
 sky130_fd_sc_hd__o21ai_0 _19059_ (.A1(_10984_),
    .A2(_13128_),
    .B1(_13129_),
    .Y(_00462_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_623 ();
 sky130_fd_sc_hd__nor2_1 _19062_ (.A(net3687),
    .B(_13078_),
    .Y(_13132_));
 sky130_fd_sc_hd__a21oi_1 _19063_ (.A1(net3503),
    .A2(_13078_),
    .B1(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__nand2_1 _19064_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .B(_13081_),
    .Y(_13134_));
 sky130_fd_sc_hd__o21ai_0 _19065_ (.A1(_13081_),
    .A2(_13133_),
    .B1(_13134_),
    .Y(_00463_));
 sky130_fd_sc_hd__nor2_1 _19066_ (.A(_09903_),
    .B(_13078_),
    .Y(_13135_));
 sky130_fd_sc_hd__a21oi_1 _19067_ (.A1(net164),
    .A2(_13078_),
    .B1(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__nand2_1 _19068_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .B(_13081_),
    .Y(_13137_));
 sky130_fd_sc_hd__o21ai_0 _19069_ (.A1(_10984_),
    .A2(_13136_),
    .B1(_13137_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_1 _19070_ (.A(_09983_),
    .B(_13078_),
    .Y(_13138_));
 sky130_fd_sc_hd__a21oi_1 _19071_ (.A1(net272),
    .A2(_13078_),
    .B1(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__nand2_1 _19072_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .B(_13081_),
    .Y(_13140_));
 sky130_fd_sc_hd__o21ai_0 _19073_ (.A1(_13081_),
    .A2(_13139_),
    .B1(_13140_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _19074_ (.A(net3495),
    .B(_13078_),
    .Y(_13141_));
 sky130_fd_sc_hd__o21ai_0 _19075_ (.A1(_10088_),
    .A2(_13078_),
    .B1(_13141_),
    .Y(_13142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_622 ();
 sky130_fd_sc_hd__mux2_1 _19077_ (.A0(_13142_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .S(_10984_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_1 _19078_ (.A(net3682),
    .B(_13078_),
    .Y(_13144_));
 sky130_fd_sc_hd__a21oi_1 _19079_ (.A1(net167),
    .A2(_13078_),
    .B1(_13144_),
    .Y(_13145_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .B(_13081_),
    .Y(_13146_));
 sky130_fd_sc_hd__o21ai_0 _19081_ (.A1(_10984_),
    .A2(_13145_),
    .B1(_13146_),
    .Y(_00467_));
 sky130_fd_sc_hd__nor2_1 _19082_ (.A(net3681),
    .B(_13078_),
    .Y(_13147_));
 sky130_fd_sc_hd__a21oi_1 _19083_ (.A1(net168),
    .A2(_13078_),
    .B1(_13147_),
    .Y(_13148_));
 sky130_fd_sc_hd__nand2_1 _19084_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B(_13081_),
    .Y(_13149_));
 sky130_fd_sc_hd__o21ai_0 _19085_ (.A1(_10984_),
    .A2(_13148_),
    .B1(_13149_),
    .Y(_00468_));
 sky130_fd_sc_hd__nor2_1 _19086_ (.A(net3679),
    .B(_13078_),
    .Y(_13150_));
 sky130_fd_sc_hd__a21oi_1 _19087_ (.A1(net169),
    .A2(_13078_),
    .B1(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand2_1 _19088_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B(_13081_),
    .Y(_13152_));
 sky130_fd_sc_hd__o21ai_0 _19089_ (.A1(_10984_),
    .A2(_13151_),
    .B1(_13152_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _19090_ (.A(net292),
    .B(_13078_),
    .Y(_13153_));
 sky130_fd_sc_hd__o21ai_0 _19091_ (.A1(net3676),
    .A2(_13078_),
    .B1(_13153_),
    .Y(_13154_));
 sky130_fd_sc_hd__mux2_1 _19092_ (.A0(_13154_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .S(_10984_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2i_1 _19093_ (.A0(net393),
    .A1(net171),
    .S(_13078_),
    .Y(_13155_));
 sky130_fd_sc_hd__nand2_1 _19094_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .B(_13081_),
    .Y(_13156_));
 sky130_fd_sc_hd__o21ai_0 _19095_ (.A1(_10984_),
    .A2(_13155_),
    .B1(_13156_),
    .Y(_00471_));
 sky130_fd_sc_hd__nor2_1 _19096_ (.A(net3674),
    .B(_13078_),
    .Y(_13157_));
 sky130_fd_sc_hd__a21oi_1 _19097_ (.A1(net481),
    .A2(_13078_),
    .B1(_13157_),
    .Y(_13158_));
 sky130_fd_sc_hd__nand2_1 _19098_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .B(_13081_),
    .Y(_13159_));
 sky130_fd_sc_hd__o21ai_0 _19099_ (.A1(_10984_),
    .A2(_13158_),
    .B1(_13159_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor3_2 _19100_ (.A(net3737),
    .B(net173),
    .C(_13076_),
    .Y(_13160_));
 sky130_fd_sc_hd__nand2_1 _19101_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B(_13081_),
    .Y(_13161_));
 sky130_fd_sc_hd__o31ai_1 _19102_ (.A1(net3675),
    .A2(_10984_),
    .A3(_13160_),
    .B1(_13161_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _19103_ (.A(net3717),
    .B(_13098_),
    .Y(_13162_));
 sky130_fd_sc_hd__o21ai_1 _19104_ (.A1(net3534),
    .A2(_13098_),
    .B1(_13162_),
    .Y(_13163_));
 sky130_fd_sc_hd__mux2_1 _19105_ (.A0(_13163_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .S(_10984_),
    .X(_00474_));
 sky130_fd_sc_hd__a21oi_1 _19106_ (.A1(net3949),
    .A2(_10980_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .Y(_13164_));
 sky130_fd_sc_hd__nor2_1 _19107_ (.A(net3708),
    .B(_13078_),
    .Y(_13165_));
 sky130_fd_sc_hd__a211oi_1 _19108_ (.A1(net3536),
    .A2(_13078_),
    .B1(_13165_),
    .C1(_13081_),
    .Y(_13166_));
 sky130_fd_sc_hd__nor2_1 _19109_ (.A(_13164_),
    .B(_13166_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _19110_ (.A(net376),
    .B(_13078_),
    .Y(_13167_));
 sky130_fd_sc_hd__a21oi_1 _19111_ (.A1(net3537),
    .A2(_13078_),
    .B1(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__nand2_1 _19112_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .B(_13081_),
    .Y(_13169_));
 sky130_fd_sc_hd__o21ai_0 _19113_ (.A1(_10984_),
    .A2(_13168_),
    .B1(_13169_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _19114_ (.A(net3724),
    .B(_13078_),
    .Y(_13170_));
 sky130_fd_sc_hd__a21oi_1 _19115_ (.A1(net177),
    .A2(net3672),
    .B1(_13170_),
    .Y(_13171_));
 sky130_fd_sc_hd__nand2_1 _19116_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .B(_13081_),
    .Y(_13172_));
 sky130_fd_sc_hd__o21ai_0 _19117_ (.A1(_10984_),
    .A2(_13171_),
    .B1(_13172_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _19118_ (.A(net403),
    .B(net3672),
    .Y(_13173_));
 sky130_fd_sc_hd__a21oi_1 _19119_ (.A1(net3530),
    .A2(net3672),
    .B1(_13173_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_1 _19120_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .B(_13081_),
    .Y(_13175_));
 sky130_fd_sc_hd__o21ai_0 _19121_ (.A1(_10984_),
    .A2(_13174_),
    .B1(_13175_),
    .Y(_00478_));
 sky130_fd_sc_hd__mux2i_1 _19122_ (.A0(net3704),
    .A1(net3519),
    .S(net3672),
    .Y(_13176_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .B(_13081_),
    .Y(_13177_));
 sky130_fd_sc_hd__o21ai_0 _19124_ (.A1(_10984_),
    .A2(_13176_),
    .B1(_13177_),
    .Y(_00479_));
 sky130_fd_sc_hd__nor2_1 _19125_ (.A(net3705),
    .B(net3672),
    .Y(_13178_));
 sky130_fd_sc_hd__a21oi_1 _19126_ (.A1(net3520),
    .A2(net3672),
    .B1(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand2_1 _19127_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .B(_13081_),
    .Y(_13180_));
 sky130_fd_sc_hd__o21ai_0 _19128_ (.A1(_10984_),
    .A2(_13179_),
    .B1(_13180_),
    .Y(_00480_));
 sky130_fd_sc_hd__maj3_4 _19129_ (.A(_10422_),
    .B(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .C(net173),
    .X(_13181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_620 ();
 sky130_fd_sc_hd__nand2_8 _19132_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .B(_10683_),
    .Y(_13184_));
 sky130_fd_sc_hd__nor3_1 _19133_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13181_),
    .C(_13184_),
    .Y(_13185_));
 sky130_fd_sc_hd__a21oi_1 _19134_ (.A1(_13071_),
    .A2(_13185_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .Y(_13186_));
 sky130_fd_sc_hd__nor2_4 _19135_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .B(_10984_),
    .Y(_13187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_619 ();
 sky130_fd_sc_hd__nor2_1 _19137_ (.A(_13186_),
    .B(_13187_),
    .Y(_00481_));
 sky130_fd_sc_hd__nor2_4 _19138_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13181_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand2_2 _19139_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__nor2_4 _19140_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13190_),
    .Y(_13191_));
 sky130_fd_sc_hd__nand2b_4 _19141_ (.A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_13192_));
 sky130_fd_sc_hd__nor2_4 _19142_ (.A(_13192_),
    .B(_13184_),
    .Y(_13193_));
 sky130_fd_sc_hd__a21oi_1 _19143_ (.A1(_13191_),
    .A2(_13193_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .Y(_13194_));
 sky130_fd_sc_hd__nor2_1 _19144_ (.A(_13187_),
    .B(_13194_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_4 _19145_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_13195_));
 sky130_fd_sc_hd__nor2_4 _19146_ (.A(_13184_),
    .B(_13195_),
    .Y(_13196_));
 sky130_fd_sc_hd__a21oi_1 _19147_ (.A1(_13191_),
    .A2(_13196_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .Y(_13197_));
 sky130_fd_sc_hd__nor2_1 _19148_ (.A(_13187_),
    .B(_13197_),
    .Y(_00483_));
 sky130_fd_sc_hd__nor2_2 _19149_ (.A(_07862_),
    .B(_10679_),
    .Y(_13198_));
 sky130_fd_sc_hd__and2_4 _19150_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_13189_),
    .X(_13199_));
 sky130_fd_sc_hd__a31oi_1 _19151_ (.A1(_13063_),
    .A2(_13198_),
    .A3(_13199_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .Y(_13200_));
 sky130_fd_sc_hd__nor2_1 _19152_ (.A(_13187_),
    .B(_13200_),
    .Y(_00484_));
 sky130_fd_sc_hd__and3_4 _19153_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_13189_),
    .X(_13201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_618 ();
 sky130_fd_sc_hd__nor2_4 _19155_ (.A(_10674_),
    .B(_13184_),
    .Y(_13203_));
 sky130_fd_sc_hd__a21oi_1 _19156_ (.A1(_13201_),
    .A2(_13203_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .Y(_13204_));
 sky130_fd_sc_hd__nor2_1 _19157_ (.A(_13187_),
    .B(_13204_),
    .Y(_00485_));
 sky130_fd_sc_hd__a21oi_1 _19158_ (.A1(_13193_),
    .A2(_13201_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .Y(_13205_));
 sky130_fd_sc_hd__nor2_1 _19159_ (.A(_13187_),
    .B(_13205_),
    .Y(_00486_));
 sky130_fd_sc_hd__a21oi_1 _19160_ (.A1(_13196_),
    .A2(_13201_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .Y(_13206_));
 sky130_fd_sc_hd__nor2_1 _19161_ (.A(_13187_),
    .B(_13206_),
    .Y(_00487_));
 sky130_fd_sc_hd__inv_1 _19162_ (.A(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .Y(_13207_));
 sky130_fd_sc_hd__maj3_4 _19163_ (.A(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B(_13207_),
    .C(net3471),
    .X(_13208_));
 sky130_fd_sc_hd__nand2_2 _19164_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13208_),
    .Y(_13209_));
 sky130_fd_sc_hd__nor2_1 _19165_ (.A(_13184_),
    .B(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__a21oi_1 _19166_ (.A1(_13071_),
    .A2(_13210_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .Y(_13211_));
 sky130_fd_sc_hd__nor2_1 _19167_ (.A(_13187_),
    .B(_13211_),
    .Y(_00488_));
 sky130_fd_sc_hd__a21oi_1 _19168_ (.A1(_10675_),
    .A2(_13210_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .Y(_13212_));
 sky130_fd_sc_hd__nor2_1 _19169_ (.A(_13187_),
    .B(_13212_),
    .Y(_00489_));
 sky130_fd_sc_hd__nor3_2 _19170_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_13209_),
    .Y(_13213_));
 sky130_fd_sc_hd__a21oi_1 _19171_ (.A1(_13193_),
    .A2(_13213_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .Y(_13214_));
 sky130_fd_sc_hd__nor2_1 _19172_ (.A(_13187_),
    .B(_13214_),
    .Y(_00490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_617 ();
 sky130_fd_sc_hd__a21oi_1 _19174_ (.A1(_13196_),
    .A2(_13213_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .Y(_13216_));
 sky130_fd_sc_hd__nor2_1 _19175_ (.A(_13187_),
    .B(_13216_),
    .Y(_00491_));
 sky130_fd_sc_hd__a21oi_1 _19176_ (.A1(_10675_),
    .A2(_13185_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .Y(_13217_));
 sky130_fd_sc_hd__nor2_1 _19177_ (.A(_13187_),
    .B(_13217_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_2 _19178_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13062_),
    .Y(_13218_));
 sky130_fd_sc_hd__nor2_2 _19179_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_13218_),
    .Y(_13219_));
 sky130_fd_sc_hd__a21oi_1 _19180_ (.A1(_13210_),
    .A2(_13219_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .Y(_13220_));
 sky130_fd_sc_hd__nor2_1 _19181_ (.A(_13187_),
    .B(_13220_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2b_4 _19182_ (.A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13221_));
 sky130_fd_sc_hd__nor2_2 _19183_ (.A(_13209_),
    .B(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__a21oi_1 _19184_ (.A1(_13203_),
    .A2(_13222_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .Y(_13223_));
 sky130_fd_sc_hd__nor2_1 _19185_ (.A(_13187_),
    .B(_13223_),
    .Y(_00494_));
 sky130_fd_sc_hd__a21oi_1 _19186_ (.A1(_13193_),
    .A2(_13222_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .Y(_13224_));
 sky130_fd_sc_hd__nor2_1 _19187_ (.A(_13187_),
    .B(_13224_),
    .Y(_00495_));
 sky130_fd_sc_hd__a21oi_1 _19188_ (.A1(_13196_),
    .A2(_13222_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .Y(_13225_));
 sky130_fd_sc_hd__nor2_1 _19189_ (.A(_13187_),
    .B(_13225_),
    .Y(_00496_));
 sky130_fd_sc_hd__and3_4 _19190_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .C(_13208_),
    .X(_13226_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_616 ();
 sky130_fd_sc_hd__a31oi_1 _19192_ (.A1(_13067_),
    .A2(_13198_),
    .A3(_13226_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .Y(_13228_));
 sky130_fd_sc_hd__nor2_1 _19193_ (.A(_13187_),
    .B(_13228_),
    .Y(_00497_));
 sky130_fd_sc_hd__and2_4 _19194_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13208_),
    .X(_13229_));
 sky130_fd_sc_hd__nand2_2 _19195_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_13229_),
    .Y(_13230_));
 sky130_fd_sc_hd__nor2_2 _19196_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__a21oi_1 _19197_ (.A1(_13203_),
    .A2(_13231_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .Y(_13232_));
 sky130_fd_sc_hd__nor2_1 _19198_ (.A(_13187_),
    .B(_13232_),
    .Y(_00498_));
 sky130_fd_sc_hd__a21oi_1 _19199_ (.A1(_13193_),
    .A2(_13231_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .Y(_13233_));
 sky130_fd_sc_hd__nor2_1 _19200_ (.A(_13187_),
    .B(_13233_),
    .Y(_00499_));
 sky130_fd_sc_hd__a21oi_1 _19201_ (.A1(_13196_),
    .A2(_13231_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .Y(_13234_));
 sky130_fd_sc_hd__nor2_1 _19202_ (.A(_13187_),
    .B(_13234_),
    .Y(_00500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_615 ();
 sky130_fd_sc_hd__a31oi_1 _19204_ (.A1(_13063_),
    .A2(_13198_),
    .A3(_13226_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .Y(_13236_));
 sky130_fd_sc_hd__nor2_1 _19205_ (.A(_13187_),
    .B(_13236_),
    .Y(_00501_));
 sky130_fd_sc_hd__and2_4 _19206_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13226_),
    .X(_13237_));
 sky130_fd_sc_hd__a21oi_1 _19207_ (.A1(_13203_),
    .A2(_13237_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .Y(_13238_));
 sky130_fd_sc_hd__nor2_1 _19208_ (.A(_13187_),
    .B(_13238_),
    .Y(_00502_));
 sky130_fd_sc_hd__nor2_1 _19209_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13239_));
 sky130_fd_sc_hd__nand2_1 _19210_ (.A(_13239_),
    .B(_13189_),
    .Y(_13240_));
 sky130_fd_sc_hd__o21ai_0 _19211_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .A2(_13081_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .Y(_13241_));
 sky130_fd_sc_hd__o31ai_1 _19212_ (.A1(_13192_),
    .A2(_13184_),
    .A3(_13240_),
    .B1(_13241_),
    .Y(_00503_));
 sky130_fd_sc_hd__a21oi_1 _19213_ (.A1(_13193_),
    .A2(_13237_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .Y(_13242_));
 sky130_fd_sc_hd__nor2_1 _19214_ (.A(_13187_),
    .B(_13242_),
    .Y(_00504_));
 sky130_fd_sc_hd__a21oi_1 _19215_ (.A1(_13196_),
    .A2(_13237_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .Y(_13243_));
 sky130_fd_sc_hd__nor2_1 _19216_ (.A(_13187_),
    .B(_13243_),
    .Y(_00505_));
 sky130_fd_sc_hd__a31oi_1 _19217_ (.A1(_13239_),
    .A2(_13189_),
    .A3(_13196_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .Y(_13244_));
 sky130_fd_sc_hd__nor2_1 _19218_ (.A(_13187_),
    .B(_13244_),
    .Y(_00506_));
 sky130_fd_sc_hd__a21oi_1 _19219_ (.A1(_13185_),
    .A2(_13219_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _19220_ (.A(_13187_),
    .B(_01645_),
    .Y(_00507_));
 sky130_fd_sc_hd__nor3_2 _19221_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13181_),
    .C(_13221_),
    .Y(_01646_));
 sky130_fd_sc_hd__a21oi_1 _19222_ (.A1(_13203_),
    .A2(_01646_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _19223_ (.A(_13187_),
    .B(_01647_),
    .Y(_00508_));
 sky130_fd_sc_hd__a21oi_1 _19224_ (.A1(_13193_),
    .A2(_01646_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _19225_ (.A(_13187_),
    .B(_01648_),
    .Y(_00509_));
 sky130_fd_sc_hd__a21oi_1 _19226_ (.A1(_13196_),
    .A2(_01646_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _19227_ (.A(_13187_),
    .B(_01649_),
    .Y(_00510_));
 sky130_fd_sc_hd__a31oi_1 _19228_ (.A1(_13067_),
    .A2(_13198_),
    .A3(_13199_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _19229_ (.A(_13187_),
    .B(_01650_),
    .Y(_00511_));
 sky130_fd_sc_hd__a21oi_1 _19230_ (.A1(_13191_),
    .A2(_13203_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .Y(_01651_));
 sky130_fd_sc_hd__nor2_1 _19231_ (.A(_13187_),
    .B(_01651_),
    .Y(_00512_));
 sky130_fd_sc_hd__or2_0 _19232_ (.A(fetch_enable_q),
    .B(net61),
    .X(_00513_));
 sky130_fd_sc_hd__a22oi_1 _19233_ (.A1(_07886_),
    .A2(_08045_),
    .B1(_08046_),
    .B2(net3834),
    .Y(_01652_));
 sky130_fd_sc_hd__o21ai_2 _19234_ (.A1(_08048_),
    .A2(_01652_),
    .B1(_08501_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_2 _19235_ (.A(_10924_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_4 _19236_ (.A(_11890_),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_609 ();
 sky130_fd_sc_hd__mux2_1 _19243_ (.A0(net57),
    .A1(net34),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_01662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_608 ();
 sky130_fd_sc_hd__mux2i_1 _19245_ (.A0(net43),
    .A1(net27),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _19246_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_607 ();
 sky130_fd_sc_hd__o211ai_1 _19248_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_01662_),
    .B1(_01665_),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_01667_));
 sky130_fd_sc_hd__mux4_2 _19249_ (.A0(net56),
    .A1(net42),
    .A2(net33),
    .A3(net51),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_01668_));
 sky130_fd_sc_hd__nand3_4 _19250_ (.A(\load_store_unit_i.data_type_q[1] ),
    .B(\load_store_unit_i.data_sign_ext_q ),
    .C(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_4 _19251_ (.A(\load_store_unit_i.data_type_q[2] ),
    .B(\load_store_unit_i.data_type_q[1] ),
    .Y(_01670_));
 sky130_fd_sc_hd__mux4_2 _19252_ (.A0(net57),
    .A1(\load_store_unit_i.rdata_q[8] ),
    .A2(\load_store_unit_i.rdata_q[16] ),
    .A3(net27),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_01671_));
 sky130_fd_sc_hd__nand2_1 _19253_ (.A(_01670_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand3_2 _19254_ (.A(_01667_),
    .B(_01669_),
    .C(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_604 ();
 sky130_fd_sc_hd__nor2_4 _19258_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Y(_01677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_603 ();
 sky130_fd_sc_hd__nor3_4 _19260_ (.A(_09572_),
    .B(net406),
    .C(_01677_),
    .Y(_01679_));
 sky130_fd_sc_hd__a21oi_4 _19261_ (.A1(net3716),
    .A2(_01677_),
    .B1(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__or2_4 _19262_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .X(_01681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_602 ();
 sky130_fd_sc_hd__mux2i_4 _19264_ (.A0(net3719),
    .A1(_09564_),
    .S(_01681_),
    .Y(_01683_));
 sky130_fd_sc_hd__nor2_1 _19265_ (.A(_01680_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__or2_4 _19266_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .X(_01685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_601 ();
 sky130_fd_sc_hd__nand4bb_4 _19268_ (.A_N(_09634_),
    .B_N(_09642_),
    .C(_09651_),
    .D(_01685_),
    .Y(_01687_));
 sky130_fd_sc_hd__a211o_4 _19269_ (.A1(_08424_),
    .A2(_08427_),
    .B1(_01685_),
    .C1(net382),
    .X(_01688_));
 sky130_fd_sc_hd__and2_4 _19270_ (.A(_01687_),
    .B(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2i_4 _19271_ (.A0(net3707),
    .A1(_09785_),
    .S(_01681_),
    .Y(_01690_));
 sky130_fd_sc_hd__nor2_2 _19272_ (.A(_01689_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_600 ();
 sky130_fd_sc_hd__mux2_8 _19274_ (.A0(_08703_),
    .A1(_09760_),
    .S(_01685_),
    .X(_01693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_599 ();
 sky130_fd_sc_hd__mux2i_4 _19276_ (.A0(net302),
    .A1(_09620_),
    .S(_01681_),
    .Y(_01695_));
 sky130_fd_sc_hd__nor2_1 _19277_ (.A(_01693_),
    .B(net447),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor3_1 _19278_ (.A(_01684_),
    .B(_01691_),
    .C(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__o311a_4 _19279_ (.A1(net3846),
    .A2(_09407_),
    .A3(_09413_),
    .B1(_09423_),
    .C1(_01681_),
    .X(_01698_));
 sky130_fd_sc_hd__a311oi_4 _19280_ (.A1(_07958_),
    .A2(_08643_),
    .A3(_08649_),
    .B1(_01681_),
    .C1(net301),
    .Y(_01699_));
 sky130_fd_sc_hd__or2_4 _19281_ (.A(_01698_),
    .B(net443),
    .X(_01700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_597 ();
 sky130_fd_sc_hd__and4_4 _19284_ (.A(_08260_),
    .B(_08281_),
    .C(_08301_),
    .D(net3761),
    .X(_01703_));
 sky130_fd_sc_hd__o211a_4 _19285_ (.A1(_09573_),
    .A2(_09711_),
    .B1(_09720_),
    .C1(_01685_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_4 _19286_ (.A(_01703_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_596 ();
 sky130_fd_sc_hd__nor2_2 _19288_ (.A(_01700_),
    .B(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__nor2_4 _19289_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .Y(_01708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_595 ();
 sky130_fd_sc_hd__a311oi_4 _19291_ (.A1(_07958_),
    .A2(_09472_),
    .A3(_09478_),
    .B1(_01708_),
    .C1(_09488_),
    .Y(_01710_));
 sky130_fd_sc_hd__a21o_4 _19292_ (.A1(net432),
    .A2(net3757),
    .B1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_594 ();
 sky130_fd_sc_hd__mux2_8 _19294_ (.A0(_08167_),
    .A1(net373),
    .S(net3758),
    .X(_01713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_591 ();
 sky130_fd_sc_hd__mux2_1 _19298_ (.A0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .S(_10740_),
    .X(_01717_));
 sky130_fd_sc_hd__a22oi_2 _19299_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_01681_),
    .B1(_01717_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_01718_));
 sky130_fd_sc_hd__o21a_1 _19300_ (.A1(_01711_),
    .A2(_01713_),
    .B1(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__nor3_1 _19301_ (.A(_01711_),
    .B(_01718_),
    .C(_01713_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _19302_ (.A(_01719_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__xnor2_1 _19303_ (.A(_01707_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nor2_1 _19304_ (.A(_01705_),
    .B(_01711_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_2 _19305_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .Y(_01724_));
 sky130_fd_sc_hd__a31oi_1 _19306_ (.A1(_08075_),
    .A2(net3820),
    .A3(net3819),
    .B1(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__a41o_4 _19307_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A3(_08028_),
    .A4(_10745_),
    .B1(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__nand2_1 _19308_ (.A(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B(_01681_),
    .Y(_01727_));
 sky130_fd_sc_hd__o21ai_4 _19309_ (.A1(_08028_),
    .A2(_01724_),
    .B1(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_589 ();
 sky130_fd_sc_hd__nor2_4 _19312_ (.A(_01726_),
    .B(_01728_),
    .Y(_01731_));
 sky130_fd_sc_hd__nor3_1 _19313_ (.A(_01705_),
    .B(_01711_),
    .C(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_2 _19314_ (.A(_01700_),
    .B(_01693_),
    .Y(_01733_));
 sky130_fd_sc_hd__o32ai_1 _19315_ (.A1(net3608),
    .A2(_01726_),
    .A3(_01728_),
    .B1(_01732_),
    .B2(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__maj3_1 _19316_ (.A(_01697_),
    .B(_01722_),
    .C(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__o21ai_0 _19317_ (.A1(_01711_),
    .A2(_01713_),
    .B1(_01718_),
    .Y(_01736_));
 sky130_fd_sc_hd__a21oi_2 _19318_ (.A1(_01707_),
    .A2(_01736_),
    .B1(_01720_),
    .Y(_01737_));
 sky130_fd_sc_hd__inv_16 _19319_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_01738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_588 ();
 sky130_fd_sc_hd__mux2i_1 _19321_ (.A0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .S(_10740_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _19322_ (.A(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B(net3759),
    .Y(_01741_));
 sky130_fd_sc_hd__o21ai_4 _19323_ (.A1(_01738_),
    .A2(_01740_),
    .B1(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__a221oi_4 _19324_ (.A1(_08786_),
    .A2(_08789_),
    .B1(_08794_),
    .B2(_08797_),
    .C1(_01685_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor4_4 _19325_ (.A(_09896_),
    .B(_09899_),
    .C(_09902_),
    .D(net3761),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_4 _19326_ (.A(_01743_),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _19327_ (.A(_01711_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _19328_ (.A(_01700_),
    .B(_01713_),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor3_1 _19329_ (.A(_01742_),
    .B(_01746_),
    .C(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__nor2_1 _19330_ (.A(_01705_),
    .B(net447),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _19331_ (.A(net397),
    .B(_01690_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _19332_ (.A(_01693_),
    .B(_01683_),
    .Y(_01751_));
 sky130_fd_sc_hd__xnor3_1 _19333_ (.A(_01749_),
    .B(_01750_),
    .C(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__xnor2_1 _19334_ (.A(_01748_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__xnor2_1 _19335_ (.A(_01737_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__maj3_4 _19336_ (.A(_01684_),
    .B(_01691_),
    .C(_01696_),
    .X(_01755_));
 sky130_fd_sc_hd__o311ai_4 _19337_ (.A1(net3846),
    .A2(_08217_),
    .A3(_08224_),
    .B1(net281),
    .C1(_01708_),
    .Y(_01756_));
 sky130_fd_sc_hd__o21a_4 _19338_ (.A1(net3691),
    .A2(_01708_),
    .B1(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2i_2 _19339_ (.A0(net3713),
    .A1(net331),
    .S(_01685_),
    .Y(_01758_));
 sky130_fd_sc_hd__mux2i_4 _19340_ (.A0(net282),
    .A1(_09863_),
    .S(_01681_),
    .Y(_01759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_587 ();
 sky130_fd_sc_hd__nor2_2 _19342_ (.A(net3648),
    .B(_01759_),
    .Y(_01761_));
 sky130_fd_sc_hd__mux2_8 _19343_ (.A0(net3711),
    .A1(net310),
    .S(net3758),
    .X(_01762_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_586 ();
 sky130_fd_sc_hd__o311ai_4 _19345_ (.A1(net3846),
    .A2(_08759_),
    .A3(_08765_),
    .B1(_08776_),
    .C1(_01708_),
    .Y(_01764_));
 sky130_fd_sc_hd__o21ai_4 _19346_ (.A1(_09935_),
    .A2(_01708_),
    .B1(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_585 ();
 sky130_fd_sc_hd__nor2_4 _19348_ (.A(_01762_),
    .B(_01765_),
    .Y(_01767_));
 sky130_fd_sc_hd__xor2_1 _19349_ (.A(_01761_),
    .B(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_583 ();
 sky130_fd_sc_hd__mux2i_4 _19352_ (.A0(net3711),
    .A1(net310),
    .S(net3758),
    .Y(_01771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_582 ();
 sky130_fd_sc_hd__nor3_1 _19354_ (.A(net3648),
    .B(_01771_),
    .C(_01759_),
    .Y(_01773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_581 ();
 sky130_fd_sc_hd__o21ai_4 _19356_ (.A1(net3691),
    .A2(_01708_),
    .B1(_01756_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_2 _19357_ (.A(_01689_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__o21ai_0 _19358_ (.A1(_01767_),
    .A2(_01773_),
    .B1(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__mux2_8 _19359_ (.A0(net3714),
    .A1(net331),
    .S(net3758),
    .X(_01778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_580 ();
 sky130_fd_sc_hd__mux2_8 _19361_ (.A0(net3727),
    .A1(_09863_),
    .S(_01681_),
    .X(_01780_));
 sky130_fd_sc_hd__a21oi_1 _19362_ (.A1(_01778_),
    .A2(_01780_),
    .B1(_01771_),
    .Y(_01781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_579 ();
 sky130_fd_sc_hd__o21a_4 _19364_ (.A1(_09935_),
    .A2(_01708_),
    .B1(_01764_),
    .X(_01783_));
 sky130_fd_sc_hd__nor3_1 _19365_ (.A(net3641),
    .B(_01762_),
    .C(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_578 ();
 sky130_fd_sc_hd__o21ai_0 _19367_ (.A1(_01781_),
    .A2(_01784_),
    .B1(_01689_),
    .Y(_01786_));
 sky130_fd_sc_hd__o211ai_1 _19368_ (.A1(_01757_),
    .A2(_01768_),
    .B1(_01777_),
    .C1(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__xor2_1 _19369_ (.A(_01755_),
    .B(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__xnor2_1 _19370_ (.A(_01754_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__xor2_1 _19371_ (.A(_01735_),
    .B(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__nor2_1 _19372_ (.A(net3648),
    .B(net3643),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _19373_ (.A(_01762_),
    .B(_01759_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_2 _19374_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__a21oi_4 _19375_ (.A1(net432),
    .A2(net3757),
    .B1(net387),
    .Y(_01794_));
 sky130_fd_sc_hd__o21ai_0 _19376_ (.A1(_01726_),
    .A2(_01728_),
    .B1(_01685_),
    .Y(_01795_));
 sky130_fd_sc_hd__o21ai_0 _19377_ (.A1(_01726_),
    .A2(_01728_),
    .B1(_01677_),
    .Y(_01796_));
 sky130_fd_sc_hd__o22ai_1 _19378_ (.A1(_09760_),
    .A2(_01795_),
    .B1(_01796_),
    .B2(_08703_),
    .Y(_01797_));
 sky130_fd_sc_hd__a21boi_0 _19379_ (.A1(_09760_),
    .A2(_01731_),
    .B1_N(_01704_),
    .Y(_01798_));
 sky130_fd_sc_hd__a21boi_0 _19380_ (.A1(_08703_),
    .A2(_01731_),
    .B1_N(_01703_),
    .Y(_01799_));
 sky130_fd_sc_hd__o22ai_1 _19381_ (.A1(_01794_),
    .A2(_01797_),
    .B1(_01798_),
    .B2(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__nor4b_1 _19382_ (.A(_01700_),
    .B(_01798_),
    .C(_01799_),
    .D_N(_01797_),
    .Y(_01801_));
 sky130_fd_sc_hd__nor2_4 _19383_ (.A(_01698_),
    .B(net443),
    .Y(_01802_));
 sky130_fd_sc_hd__nor4_1 _19384_ (.A(_01802_),
    .B(_01705_),
    .C(_01711_),
    .D(_01731_),
    .Y(_01803_));
 sky130_fd_sc_hd__a211oi_1 _19385_ (.A1(_01800_),
    .A2(_01707_),
    .B1(_01801_),
    .C1(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__xnor3_1 _19386_ (.A(_01804_),
    .B(_01697_),
    .C(_01721_),
    .X(_01805_));
 sky130_fd_sc_hd__xnor3_1 _19387_ (.A(_01723_),
    .B(_01731_),
    .C(_01733_),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_1 _19388_ (.A(_01700_),
    .B(net398),
    .Y(_01807_));
 sky130_fd_sc_hd__mux2_1 _19389_ (.A0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .S(_10740_),
    .X(_01808_));
 sky130_fd_sc_hd__a22oi_2 _19390_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(net3759),
    .B1(_01808_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_01809_));
 sky130_fd_sc_hd__inv_1 _19391_ (.A(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_2 _19392_ (.A(_01711_),
    .B(_01693_),
    .Y(_01811_));
 sky130_fd_sc_hd__maj3_4 _19393_ (.A(_01807_),
    .B(_01810_),
    .C(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__xor3_1 _19394_ (.A(net3608),
    .B(_01731_),
    .C(_01733_),
    .X(_01813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_577 ();
 sky130_fd_sc_hd__a21o_4 _19396_ (.A1(net3716),
    .A2(_01677_),
    .B1(_01679_),
    .X(_01815_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(_01802_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_576 ();
 sky130_fd_sc_hd__mux2i_4 _19399_ (.A0(_08703_),
    .A1(_09760_),
    .S(_01685_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _19400_ (.A(_01794_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__maj3_1 _19401_ (.A(_01816_),
    .B(_01809_),
    .C(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__nor2_1 _19402_ (.A(_01680_),
    .B(net447),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _19403_ (.A(_01683_),
    .B(_01689_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _19404_ (.A(_01690_),
    .B(net3648),
    .Y(_01823_));
 sky130_fd_sc_hd__xnor3_1 _19405_ (.A(_01821_),
    .B(_01822_),
    .C(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__o21ai_0 _19406_ (.A1(_01813_),
    .A2(_01820_),
    .B1(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__o21ai_2 _19407_ (.A1(net3585),
    .A2(_01812_),
    .B1(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_573 ();
 sky130_fd_sc_hd__nor4_2 _19411_ (.A(_01680_),
    .B(_01683_),
    .C(_01689_),
    .D(net447),
    .Y(_01830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_572 ();
 sky130_fd_sc_hd__o22ai_2 _19413_ (.A1(_01683_),
    .A2(_01689_),
    .B1(net447),
    .B2(_01680_),
    .Y(_01832_));
 sky130_fd_sc_hd__o21ai_4 _19414_ (.A1(net3607),
    .A2(_01830_),
    .B1(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__and3_1 _19415_ (.A(_01805_),
    .B(_01826_),
    .C(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__maj3_1 _19416_ (.A(_01805_),
    .B(_01826_),
    .C(_01833_),
    .X(_01835_));
 sky130_fd_sc_hd__o21ai_2 _19417_ (.A1(_01793_),
    .A2(_01834_),
    .B1(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor4_1 _19418_ (.A(_01805_),
    .B(_01826_),
    .C(_01833_),
    .D(_01793_),
    .Y(_01837_));
 sky130_fd_sc_hd__a21oi_4 _19419_ (.A1(_01790_),
    .A2(_01836_),
    .B1(net3561),
    .Y(_01838_));
 sky130_fd_sc_hd__mux2i_1 _19420_ (.A0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .S(_10740_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _19421_ (.A(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .B(net3759),
    .Y(_01840_));
 sky130_fd_sc_hd__o21ai_4 _19422_ (.A1(_01738_),
    .A2(_01839_),
    .B1(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__a211o_4 _19423_ (.A1(_08927_),
    .A2(_08930_),
    .B1(_08938_),
    .C1(_01685_),
    .X(_01842_));
 sky130_fd_sc_hd__o31a_1 _19424_ (.A1(_09961_),
    .A2(_09982_),
    .A3(net3761),
    .B1(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__nor2_1 _19425_ (.A(_01711_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _19426_ (.A(_01700_),
    .B(_01745_),
    .Y(_01845_));
 sky130_fd_sc_hd__xnor3_1 _19427_ (.A(_01841_),
    .B(_01844_),
    .C(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__nor4_1 _19428_ (.A(_01700_),
    .B(net3651),
    .C(_01713_),
    .D(_01745_),
    .Y(_01847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_571 ();
 sky130_fd_sc_hd__o22ai_1 _19430_ (.A1(_01700_),
    .A2(net445),
    .B1(_01745_),
    .B2(net3651),
    .Y(_01849_));
 sky130_fd_sc_hd__o21ai_2 _19431_ (.A1(_01742_),
    .A2(_01847_),
    .B1(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _19432_ (.A(_01705_),
    .B(_01683_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_2 _19433_ (.A(net450),
    .B(net445),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_2 _19434_ (.A(_01693_),
    .B(_01690_),
    .Y(_01853_));
 sky130_fd_sc_hd__xnor3_1 _19435_ (.A(_01851_),
    .B(_01852_),
    .C(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__xor3_1 _19436_ (.A(_01846_),
    .B(_01850_),
    .C(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__maj3_1 _19437_ (.A(_01749_),
    .B(_01750_),
    .C(_01751_),
    .X(_01856_));
 sky130_fd_sc_hd__nor2_1 _19438_ (.A(net397),
    .B(_01775_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _19439_ (.A(_01689_),
    .B(_01759_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_2 _19440_ (.A(net3648),
    .B(_01765_),
    .Y(_01859_));
 sky130_fd_sc_hd__xor3_1 _19441_ (.A(_01857_),
    .B(_01858_),
    .C(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__maj3_2 _19442_ (.A(_01776_),
    .B(_01761_),
    .C(_01767_),
    .X(_01861_));
 sky130_fd_sc_hd__xnor3_1 _19443_ (.A(_01856_),
    .B(_01860_),
    .C(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__maj3_1 _19444_ (.A(_01737_),
    .B(_01748_),
    .C(_01752_),
    .X(_01863_));
 sky130_fd_sc_hd__xnor2_1 _19445_ (.A(_01862_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__xnor2_2 _19446_ (.A(_01855_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_570 ();
 sky130_fd_sc_hd__mux2i_4 _19448_ (.A0(_08917_),
    .A1(_10010_),
    .S(net3760),
    .Y(_01867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_569 ();
 sky130_fd_sc_hd__nor2_4 _19450_ (.A(_01762_),
    .B(_01867_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_4 _19451_ (.A(_01757_),
    .B(net3645),
    .Y(_01870_));
 sky130_fd_sc_hd__nor3_2 _19452_ (.A(_01689_),
    .B(_01775_),
    .C(_01767_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor3_2 _19453_ (.A(_01762_),
    .B(net3646),
    .C(_01776_),
    .Y(_01872_));
 sky130_fd_sc_hd__nor3_1 _19454_ (.A(_01870_),
    .B(_01871_),
    .C(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__o211ai_1 _19455_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01761_),
    .C1(_01870_),
    .Y(_01874_));
 sky130_fd_sc_hd__or3_1 _19456_ (.A(_01761_),
    .B(_01871_),
    .C(_01872_),
    .X(_01875_));
 sky130_fd_sc_hd__o211ai_1 _19457_ (.A1(_01755_),
    .A2(_01873_),
    .B1(_01874_),
    .C1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__xnor2_2 _19458_ (.A(_01869_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__maj3_4 _19459_ (.A(_01735_),
    .B(_01754_),
    .C(_01788_),
    .X(_01878_));
 sky130_fd_sc_hd__xor2_1 _19460_ (.A(_01877_),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__xnor2_2 _19461_ (.A(_01865_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__xnor2_1 _19462_ (.A(_01838_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__maj3_1 _19463_ (.A(_01826_),
    .B(_01833_),
    .C(_01793_),
    .X(_01882_));
 sky130_fd_sc_hd__and3_1 _19464_ (.A(_01826_),
    .B(_01833_),
    .C(_01793_),
    .X(_01883_));
 sky130_fd_sc_hd__a211oi_1 _19465_ (.A1(_01805_),
    .A2(_01882_),
    .B1(_01883_),
    .C1(_01837_),
    .Y(_01884_));
 sky130_fd_sc_hd__xnor2_1 _19466_ (.A(_01790_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_8 _19467_ (.A(net3671),
    .B(_01688_),
    .Y(_01886_));
 sky130_fd_sc_hd__mux2_8 _19468_ (.A0(net302),
    .A1(_09620_),
    .S(_01681_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_8 _19469_ (.A0(net3719),
    .A1(_09564_),
    .S(_01681_),
    .X(_01888_));
 sky130_fd_sc_hd__a22oi_1 _19470_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01778_),
    .B2(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__mux2_8 _19471_ (.A0(net3707),
    .A1(_09785_),
    .S(_01681_),
    .X(_01890_));
 sky130_fd_sc_hd__a41oi_1 _19472_ (.A1(_01888_),
    .A2(_01886_),
    .A3(_01887_),
    .A4(_01778_),
    .B1(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__or2_4 _19473_ (.A(_01889_),
    .B(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__nand2_2 _19474_ (.A(net3585),
    .B(_01812_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor2_1 _19475_ (.A(net442),
    .B(_01758_),
    .Y(_01894_));
 sky130_fd_sc_hd__a22oi_1 _19476_ (.A1(_01821_),
    .A2(net3607),
    .B1(net3604),
    .B2(_01691_),
    .Y(_01895_));
 sky130_fd_sc_hd__a32oi_1 _19477_ (.A1(_01821_),
    .A2(_01822_),
    .A3(net3607),
    .B1(_01820_),
    .B2(_01813_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor3_1 _19478_ (.A(net3585),
    .B(_01812_),
    .C(_01833_),
    .Y(_01897_));
 sky130_fd_sc_hd__o22ai_2 _19479_ (.A1(_01893_),
    .A2(_01895_),
    .B1(_01896_),
    .B2(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _19480_ (.A(net3607),
    .B(_01832_),
    .Y(_01899_));
 sky130_fd_sc_hd__mux2_4 _19481_ (.A0(_01830_),
    .A1(_01899_),
    .S(_01893_),
    .X(_01900_));
 sky130_fd_sc_hd__xnor2_1 _19482_ (.A(_01805_),
    .B(_01793_),
    .Y(_01901_));
 sky130_fd_sc_hd__o21ai_0 _19483_ (.A1(_01898_),
    .A2(_01900_),
    .B1(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__or3_1 _19484_ (.A(_01898_),
    .B(_01900_),
    .C(_01901_),
    .X(_01903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_568 ();
 sky130_fd_sc_hd__o21ai_0 _19486_ (.A1(net3656),
    .A2(_01889_),
    .B1(net3641),
    .Y(_01905_));
 sky130_fd_sc_hd__or3_1 _19487_ (.A(net3641),
    .B(_01889_),
    .C(_01891_),
    .X(_01906_));
 sky130_fd_sc_hd__nand2_1 _19488_ (.A(_01886_),
    .B(_01887_),
    .Y(_01907_));
 sky130_fd_sc_hd__nor3_1 _19489_ (.A(net3658),
    .B(net3649),
    .C(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__a32o_1 _19490_ (.A1(net3645),
    .A2(_01905_),
    .A3(_01906_),
    .B1(_01870_),
    .B2(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_2 _19491_ (.A(_01794_),
    .B(_01815_),
    .Y(_01910_));
 sky130_fd_sc_hd__mux2_1 _19492_ (.A0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .S(_10740_),
    .X(_01911_));
 sky130_fd_sc_hd__a22oi_2 _19493_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_01681_),
    .B1(_01911_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_01912_));
 sky130_fd_sc_hd__a211oi_2 _19494_ (.A1(net3671),
    .A2(_01688_),
    .B1(_01698_),
    .C1(net443),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2b_2 _19495_ (.A_N(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2b_1 _19496_ (.A(_01913_),
    .B_N(_01912_),
    .Y(_01915_));
 sky130_fd_sc_hd__a21oi_1 _19497_ (.A1(_01910_),
    .A2(_01914_),
    .B1(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _19498_ (.A(_01690_),
    .B(_01762_),
    .Y(_01917_));
 sky130_fd_sc_hd__xnor3_1 _19499_ (.A(_01894_),
    .B(_01907_),
    .C(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__xnor3_1 _19500_ (.A(_01807_),
    .B(_01809_),
    .C(_01811_),
    .X(_01919_));
 sky130_fd_sc_hd__maj3_1 _19501_ (.A(_01916_),
    .B(_01918_),
    .C(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__xnor3_1 _19502_ (.A(_01806_),
    .B(_01812_),
    .C(_01824_),
    .X(_01921_));
 sky130_fd_sc_hd__maj3_1 _19503_ (.A(_01909_),
    .B(_01920_),
    .C(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__a21oi_1 _19504_ (.A1(_01902_),
    .A2(_01903_),
    .B1(net3572),
    .Y(_01923_));
 sky130_fd_sc_hd__nand3_1 _19505_ (.A(_01902_),
    .B(_01903_),
    .C(net3572),
    .Y(_01924_));
 sky130_fd_sc_hd__o31a_1 _19506_ (.A1(_01870_),
    .A2(_01892_),
    .A3(_01923_),
    .B1(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__nor2_4 _19507_ (.A(net3655),
    .B(_01762_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_2 _19508_ (.A(net3604),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__mux2i_1 _19509_ (.A0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .S(_10740_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _19510_ (.A(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B(_01681_),
    .Y(_01929_));
 sky130_fd_sc_hd__o21a_4 _19511_ (.A1(_01738_),
    .A2(_01928_),
    .B1(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__nand2_1 _19512_ (.A(_01794_),
    .B(_01886_),
    .Y(_01931_));
 sky130_fd_sc_hd__nand2_1 _19513_ (.A(_01802_),
    .B(_01778_),
    .Y(_01932_));
 sky130_fd_sc_hd__maj3_2 _19514_ (.A(_01930_),
    .B(_01931_),
    .C(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__xnor2_1 _19515_ (.A(_01913_),
    .B(_01912_),
    .Y(_01934_));
 sky130_fd_sc_hd__xor2_1 _19516_ (.A(_01910_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nor2_1 _19517_ (.A(net3658),
    .B(_01762_),
    .Y(_01936_));
 sky130_fd_sc_hd__a21oi_1 _19518_ (.A1(_01887_),
    .A2(_01778_),
    .B1(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__maj3_1 _19519_ (.A(_01933_),
    .B(_01935_),
    .C(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_567 ();
 sky130_fd_sc_hd__o22ai_1 _19521_ (.A1(_01700_),
    .A2(_01689_),
    .B1(_01912_),
    .B2(net398),
    .Y(_01940_));
 sky130_fd_sc_hd__nand2_1 _19522_ (.A(net398),
    .B(_01912_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand3_1 _19523_ (.A(_01811_),
    .B(_01940_),
    .C(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_566 ();
 sky130_fd_sc_hd__o211ai_1 _19525_ (.A1(net398),
    .A2(_01915_),
    .B1(_01914_),
    .C1(_01693_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _19526_ (.A(_01711_),
    .B(_01914_),
    .Y(_01945_));
 sky130_fd_sc_hd__nand3_1 _19527_ (.A(_01942_),
    .B(_01944_),
    .C(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__xnor2_1 _19528_ (.A(_01816_),
    .B(_01809_),
    .Y(_01947_));
 sky130_fd_sc_hd__xnor2_1 _19529_ (.A(_01918_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__xnor2_1 _19530_ (.A(_01946_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__a21bo_4 _19531_ (.A1(_01927_),
    .A2(_01938_),
    .B1_N(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__or3_4 _19532_ (.A(_01927_),
    .B(_01933_),
    .C(_01935_),
    .X(_01951_));
 sky130_fd_sc_hd__xnor3_1 _19533_ (.A(_01909_),
    .B(_01920_),
    .C(net3579),
    .X(_01952_));
 sky130_fd_sc_hd__a21oi_2 _19534_ (.A1(_01950_),
    .A2(_01951_),
    .B1(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__xnor3_1 _19535_ (.A(_01930_),
    .B(_01931_),
    .C(_01932_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_1 _19536_ (.A(_01887_),
    .B(_01778_),
    .Y(_01955_));
 sky130_fd_sc_hd__o21ai_2 _19537_ (.A1(_01738_),
    .A2(_01928_),
    .B1(_01929_),
    .Y(_01956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_565 ();
 sky130_fd_sc_hd__a221oi_2 _19539_ (.A1(net432),
    .A2(net3757),
    .B1(net3671),
    .B2(_01688_),
    .C1(net388),
    .Y(_01958_));
 sky130_fd_sc_hd__maj3_1 _19540_ (.A(_01802_),
    .B(_01956_),
    .C(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__o2111ai_1 _19541_ (.A1(_01956_),
    .A2(_01958_),
    .B1(_01802_),
    .C1(net3655),
    .D1(_01778_),
    .Y(_01960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_564 ();
 sky130_fd_sc_hd__o211ai_1 _19543_ (.A1(net3655),
    .A2(net3649),
    .B1(_01956_),
    .C1(_01958_),
    .Y(_01962_));
 sky130_fd_sc_hd__o211ai_1 _19544_ (.A1(_01955_),
    .A2(_01959_),
    .B1(_01960_),
    .C1(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor3_1 _19545_ (.A(_01910_),
    .B(_01936_),
    .C(_01934_),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_1 _19546_ (.A(_01963_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__mux2i_1 _19547_ (.A0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .S(_10740_),
    .Y(_01966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_563 ();
 sky130_fd_sc_hd__nand2_1 _19549_ (.A(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B(net3759),
    .Y(_01968_));
 sky130_fd_sc_hd__o21ai_4 _19550_ (.A1(_01738_),
    .A2(_01966_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_1 _19551_ (.A(_01700_),
    .B(_01762_),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _19552_ (.A(_01711_),
    .B(net3649),
    .Y(_01971_));
 sky130_fd_sc_hd__maj3_4 _19553_ (.A(_01969_),
    .B(_01970_),
    .C(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__nand2_1 _19554_ (.A(_01926_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__xnor2_1 _19555_ (.A(_01700_),
    .B(_01969_),
    .Y(_01974_));
 sky130_fd_sc_hd__xnor2_1 _19556_ (.A(net3649),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_562 ();
 sky130_fd_sc_hd__mux2i_1 _19558_ (.A0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .S(_10740_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand2_1 _19559_ (.A(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B(net3759),
    .Y(_01978_));
 sky130_fd_sc_hd__o21ai_4 _19560_ (.A1(_01738_),
    .A2(_01977_),
    .B1(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__and3_4 _19561_ (.A(net3640),
    .B(net3645),
    .C(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_2 _19562_ (.A(_01975_),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a21oi_1 _19563_ (.A1(_01965_),
    .A2(_01973_),
    .B1(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__o211ai_1 _19564_ (.A1(_01926_),
    .A2(_01972_),
    .B1(_01975_),
    .C1(_01980_),
    .Y(_01983_));
 sky130_fd_sc_hd__o21ai_0 _19565_ (.A1(_01926_),
    .A2(_01972_),
    .B1(_01954_),
    .Y(_01984_));
 sky130_fd_sc_hd__a31oi_1 _19566_ (.A1(_01973_),
    .A2(_01983_),
    .A3(_01984_),
    .B1(_01965_),
    .Y(_01985_));
 sky130_fd_sc_hd__a21oi_2 _19567_ (.A1(_01954_),
    .A2(_01982_),
    .B1(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__a21o_1 _19568_ (.A1(_01927_),
    .A2(_01935_),
    .B1(_01937_),
    .X(_01987_));
 sky130_fd_sc_hd__nor3_1 _19569_ (.A(_01927_),
    .B(_01933_),
    .C(_01935_),
    .Y(_01988_));
 sky130_fd_sc_hd__a221oi_1 _19570_ (.A1(_01935_),
    .A2(_01937_),
    .B1(_01987_),
    .B2(_01933_),
    .C1(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__xnor2_1 _19571_ (.A(_01949_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__a311oi_2 _19572_ (.A1(_01952_),
    .A2(_01950_),
    .A3(_01951_),
    .B1(_01986_),
    .C1(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _19573_ (.A(_01898_),
    .B(_01900_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _19574_ (.A(_01870_),
    .B(_01892_),
    .Y(_01993_));
 sky130_fd_sc_hd__xnor2_1 _19575_ (.A(_01993_),
    .B(_01922_),
    .Y(_01994_));
 sky130_fd_sc_hd__xor3_1 _19576_ (.A(_01992_),
    .B(_01901_),
    .C(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__o21ai_2 _19577_ (.A1(_01953_),
    .A2(_01991_),
    .B1(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__maj3_4 _19578_ (.A(_01885_),
    .B(_01925_),
    .C(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__xor2_4 _19579_ (.A(net3523),
    .B(net3522),
    .X(_01998_));
 sky130_fd_sc_hd__nor2_4 _19580_ (.A(net3785),
    .B(net3744),
    .Y(_01999_));
 sky130_fd_sc_hd__or3_4 _19581_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .C(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_560 ();
 sky130_fd_sc_hd__mux2i_4 _19584_ (.A0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .A1(_01998_),
    .S(_02000_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _19585_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .Y(_02004_));
 sky130_fd_sc_hd__o21ai_2 _19586_ (.A1(net3937),
    .A2(_02003_),
    .B1(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__and2_4 _19587_ (.A(net384),
    .B(_10937_),
    .X(_02006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_559 ();
 sky130_fd_sc_hd__nand2_1 _19589_ (.A(net3519),
    .B(_02006_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor3_2 _19590_ (.A(net3725),
    .B(_08050_),
    .C(net472),
    .Y(_02009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_557 ();
 sky130_fd_sc_hd__nor2_4 _19593_ (.A(net3818),
    .B(_11012_),
    .Y(_02012_));
 sky130_fd_sc_hd__xnor2_1 _19594_ (.A(_08737_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_556 ();
 sky130_fd_sc_hd__a21oi_4 _19596_ (.A1(net3622),
    .A2(_10600_),
    .B1(net3818),
    .Y(_02015_));
 sky130_fd_sc_hd__xnor2_4 _19597_ (.A(_08359_),
    .B(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_554 ();
 sky130_fd_sc_hd__nand2_1 _19600_ (.A(net3599),
    .B(net3603),
    .Y(_02019_));
 sky130_fd_sc_hd__or3_4 _19601_ (.A(net3725),
    .B(net336),
    .C(net472),
    .X(_02020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_553 ();
 sky130_fd_sc_hd__nand2_1 _19603_ (.A(_10269_),
    .B(_02020_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_2 _19604_ (.A(_02019_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_552 ();
 sky130_fd_sc_hd__nor2_1 _19606_ (.A(_10203_),
    .B(net3603),
    .Y(_02025_));
 sky130_fd_sc_hd__a21oi_1 _19607_ (.A1(net3594),
    .A2(net3603),
    .B1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _19608_ (.A(net3621),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__o21ai_1 _19609_ (.A1(net3621),
    .A2(_02023_),
    .B1(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _19610_ (.A(net3598),
    .B(net3603),
    .Y(_02029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_551 ();
 sky130_fd_sc_hd__nand2_1 _19612_ (.A(_10336_),
    .B(_02020_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _19613_ (.A(_02029_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_10452_),
    .B(_02020_),
    .Y(_02033_));
 sky130_fd_sc_hd__o21ai_1 _19615_ (.A1(net3597),
    .A2(_02020_),
    .B1(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__mux2i_1 _19616_ (.A0(_02032_),
    .A1(_02034_),
    .S(net3619),
    .Y(_02035_));
 sky130_fd_sc_hd__nand2_1 _19617_ (.A(_08031_),
    .B(net3619),
    .Y(_02036_));
 sky130_fd_sc_hd__xnor2_1 _19618_ (.A(net308),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_550 ();
 sky130_fd_sc_hd__mux2i_1 _19620_ (.A0(_02028_),
    .A1(_02035_),
    .S(net3578),
    .Y(_02039_));
 sky130_fd_sc_hd__mux2i_1 _19621_ (.A0(net3615),
    .A1(_09907_),
    .S(_02020_),
    .Y(_02040_));
 sky130_fd_sc_hd__mux2i_1 _19622_ (.A0(_08810_),
    .A1(_09986_),
    .S(_02020_),
    .Y(_02041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_549 ();
 sky130_fd_sc_hd__mux2i_1 _19624_ (.A0(_02040_),
    .A1(_02041_),
    .S(net3619),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _19625_ (.A(_10098_),
    .B(_02020_),
    .Y(_02044_));
 sky130_fd_sc_hd__o21ai_1 _19626_ (.A1(net3601),
    .A2(_02020_),
    .B1(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_1 _19627_ (.A(_10173_),
    .B(_02020_),
    .Y(_02046_));
 sky130_fd_sc_hd__o21ai_2 _19628_ (.A1(net3600),
    .A2(_02020_),
    .B1(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__mux2i_1 _19629_ (.A0(_02045_),
    .A1(_02047_),
    .S(net3619),
    .Y(_02048_));
 sky130_fd_sc_hd__mux2i_1 _19630_ (.A0(_02043_),
    .A1(_02048_),
    .S(net3578),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _19631_ (.A(net3818),
    .B(_10600_),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_2 _19632_ (.A(_10550_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_548 ();
 sky130_fd_sc_hd__mux2i_2 _19634_ (.A0(_02039_),
    .A1(_02049_),
    .S(net3558),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _19635_ (.A(_10427_),
    .B(net3603),
    .Y(_02054_));
 sky130_fd_sc_hd__a21oi_4 _19636_ (.A1(net3620),
    .A2(net3603),
    .B1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__xnor2_4 _19637_ (.A(net3623),
    .B(_02015_),
    .Y(_02056_));
 sky130_fd_sc_hd__or3b_4 _19638_ (.A(net372),
    .B(net3725),
    .C_N(net336),
    .X(_02057_));
 sky130_fd_sc_hd__nor2_4 _19639_ (.A(_10931_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21o_1 _19640_ (.A1(net3622),
    .A2(_10600_),
    .B1(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__and3_4 _19641_ (.A(_02055_),
    .B(_02056_),
    .C(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__a21oi_4 _19642_ (.A1(_02016_),
    .A2(_02053_),
    .B1(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_547 ();
 sky130_fd_sc_hd__a21oi_2 _19644_ (.A1(_02055_),
    .A2(_02058_),
    .B1(net3560),
    .Y(_02063_));
 sky130_fd_sc_hd__a21oi_2 _19645_ (.A1(net3560),
    .A2(_02061_),
    .B1(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_546 ();
 sky130_fd_sc_hd__mux2i_1 _19647_ (.A0(_02023_),
    .A1(_02032_),
    .S(net3619),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _19648_ (.A(net3619),
    .B(_02055_),
    .Y(_02067_));
 sky130_fd_sc_hd__o21ai_2 _19649_ (.A1(net3619),
    .A2(_02034_),
    .B1(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_545 ();
 sky130_fd_sc_hd__mux2i_2 _19651_ (.A0(_02066_),
    .A1(_02068_),
    .S(net3578),
    .Y(_02070_));
 sky130_fd_sc_hd__mux2i_1 _19652_ (.A0(_02041_),
    .A1(_02045_),
    .S(net3619),
    .Y(_02071_));
 sky130_fd_sc_hd__nand2_1 _19653_ (.A(net3619),
    .B(_02026_),
    .Y(_02072_));
 sky130_fd_sc_hd__o21ai_2 _19654_ (.A1(net3619),
    .A2(_02047_),
    .B1(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_544 ();
 sky130_fd_sc_hd__mux2i_2 _19656_ (.A0(_02071_),
    .A1(_02073_),
    .S(net3578),
    .Y(_02075_));
 sky130_fd_sc_hd__mux2i_2 _19657_ (.A0(_02070_),
    .A1(_02075_),
    .S(net3558),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_8 _19658_ (.A(_02055_),
    .B(_02058_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_4 _19659_ (.A(_02077_),
    .B(_02056_),
    .Y(_02078_));
 sky130_fd_sc_hd__o21ai_2 _19660_ (.A1(_02056_),
    .A2(_02076_),
    .B1(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _19661_ (.A(_09797_),
    .B(_02020_),
    .Y(_02080_));
 sky130_fd_sc_hd__o21ai_1 _19662_ (.A1(_08988_),
    .A2(_02020_),
    .B1(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__mux2i_1 _19663_ (.A0(net3592),
    .A1(_09730_),
    .S(_02020_),
    .Y(_02082_));
 sky130_fd_sc_hd__mux2i_1 _19664_ (.A0(_02081_),
    .A1(_02082_),
    .S(net3619),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _19665_ (.A(net438),
    .B(_02020_),
    .Y(_02084_));
 sky130_fd_sc_hd__o21ai_0 _19666_ (.A1(net3617),
    .A2(_02020_),
    .B1(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__mux2i_1 _19667_ (.A0(_02040_),
    .A1(_02085_),
    .S(net3621),
    .Y(_02086_));
 sky130_fd_sc_hd__mux2i_1 _19668_ (.A0(_02083_),
    .A1(_02086_),
    .S(net3578),
    .Y(_02087_));
 sky130_fd_sc_hd__mux2i_2 _19669_ (.A0(net3589),
    .A1(net3613),
    .S(_02020_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _19670_ (.A(net3590),
    .B(_02020_),
    .Y(_02089_));
 sky130_fd_sc_hd__nor2_1 _19671_ (.A(net3588),
    .B(net3603),
    .Y(_02090_));
 sky130_fd_sc_hd__or3_1 _19672_ (.A(net3619),
    .B(_02089_),
    .C(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__o21ai_1 _19673_ (.A1(net3621),
    .A2(_02088_),
    .B1(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__mux2i_1 _19674_ (.A0(net3591),
    .A1(_09663_),
    .S(_02020_),
    .Y(_02093_));
 sky130_fd_sc_hd__mux2i_1 _19675_ (.A0(_09214_),
    .A1(_09593_),
    .S(_02020_),
    .Y(_02094_));
 sky130_fd_sc_hd__mux2i_1 _19676_ (.A0(_02093_),
    .A1(_02094_),
    .S(net3619),
    .Y(_02095_));
 sky130_fd_sc_hd__mux2i_1 _19677_ (.A0(_02092_),
    .A1(_02095_),
    .S(net3578),
    .Y(_02096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_543 ();
 sky130_fd_sc_hd__mux2i_2 _19679_ (.A0(_02087_),
    .A1(_02096_),
    .S(net3558),
    .Y(_02098_));
 sky130_fd_sc_hd__mux2i_1 _19680_ (.A0(_09214_),
    .A1(_09593_),
    .S(net3603),
    .Y(_02099_));
 sky130_fd_sc_hd__mux2i_1 _19681_ (.A0(net3591),
    .A1(_09663_),
    .S(net3603),
    .Y(_02100_));
 sky130_fd_sc_hd__mux2i_1 _19682_ (.A0(_02099_),
    .A1(_02100_),
    .S(net3619),
    .Y(_02101_));
 sky130_fd_sc_hd__mux2i_2 _19683_ (.A0(net3589),
    .A1(net3613),
    .S(net3603),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _19684_ (.A(net3588),
    .B(_02020_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _19685_ (.A(net3590),
    .B(net3603),
    .Y(_02104_));
 sky130_fd_sc_hd__or3_1 _19686_ (.A(net3621),
    .B(_02103_),
    .C(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__o21ai_1 _19687_ (.A1(net3619),
    .A2(_02102_),
    .B1(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__mux2i_1 _19688_ (.A0(_02101_),
    .A1(_02106_),
    .S(net3578),
    .Y(_02107_));
 sky130_fd_sc_hd__mux2i_1 _19689_ (.A0(net3615),
    .A1(_09907_),
    .S(net3603),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _19690_ (.A(net438),
    .B(net3603),
    .Y(_02109_));
 sky130_fd_sc_hd__o21ai_1 _19691_ (.A1(net3617),
    .A2(net3603),
    .B1(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__mux2i_1 _19692_ (.A0(_02108_),
    .A1(_02110_),
    .S(net3619),
    .Y(_02111_));
 sky130_fd_sc_hd__mux2i_1 _19693_ (.A0(net3592),
    .A1(_09730_),
    .S(net3603),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _19694_ (.A(_09797_),
    .B(net3603),
    .Y(_02113_));
 sky130_fd_sc_hd__o21ai_2 _19695_ (.A1(_08988_),
    .A2(net3603),
    .B1(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__mux2i_1 _19696_ (.A0(_02112_),
    .A1(_02114_),
    .S(net3619),
    .Y(_02115_));
 sky130_fd_sc_hd__mux2i_1 _19697_ (.A0(_02111_),
    .A1(_02115_),
    .S(net3578),
    .Y(_02116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_542 ();
 sky130_fd_sc_hd__mux2_1 _19699_ (.A0(_02107_),
    .A1(_02116_),
    .S(net3558),
    .X(_02118_));
 sky130_fd_sc_hd__nand2_1 _19700_ (.A(_02016_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__o211ai_1 _19701_ (.A1(_02016_),
    .A2(_02098_),
    .B1(_02119_),
    .C1(net3560),
    .Y(_02120_));
 sky130_fd_sc_hd__o21ai_2 _19702_ (.A1(net3560),
    .A2(_02079_),
    .B1(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__nor3b_2 _19703_ (.A(net372),
    .B(net3725),
    .C_N(net384),
    .Y(_02122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_541 ();
 sky130_fd_sc_hd__nor2_4 _19705_ (.A(net372),
    .B(net335),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2b_4 _19706_ (.A_N(_10942_),
    .B(_10940_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand2_4 _19707_ (.A(_10939_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_8 _19708_ (.A(_02124_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_540 ();
 sky130_fd_sc_hd__and4_4 _19710_ (.A(net3940),
    .B(net3943),
    .C(net3936),
    .D(_08058_),
    .X(_02129_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_539 ();
 sky130_fd_sc_hd__nand2_1 _19712_ (.A(net3616),
    .B(net3615),
    .Y(_02131_));
 sky130_fd_sc_hd__xnor2_1 _19713_ (.A(_02129_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand3_4 _19714_ (.A(net3940),
    .B(_08010_),
    .C(_08058_),
    .Y(_02133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_538 ();
 sky130_fd_sc_hd__inv_2 _19716_ (.A(_02125_),
    .Y(_02135_));
 sky130_fd_sc_hd__o21ai_4 _19717_ (.A1(_10937_),
    .A2(_02135_),
    .B1(_02124_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_8 _19718_ (.A(_02133_),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_537 ();
 sky130_fd_sc_hd__o21ai_0 _19720_ (.A1(net3616),
    .A2(net3615),
    .B1(_02137_),
    .Y(_02139_));
 sky130_fd_sc_hd__a21oi_1 _19721_ (.A1(_02127_),
    .A2(_02132_),
    .B1(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__a221oi_2 _19722_ (.A1(net3603),
    .A2(_02064_),
    .B1(_02121_),
    .B2(net3602),
    .C1(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand3_2 _19723_ (.A(net3745),
    .B(_02008_),
    .C(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__o21ai_4 _19724_ (.A1(net3745),
    .A2(_02005_),
    .B1(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand3_4 _19725_ (.A(_11705_),
    .B(_01655_),
    .C(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__o21ai_4 _19726_ (.A1(net3469),
    .A2(_01673_),
    .B1(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_536 ();
 sky130_fd_sc_hd__and3_4 _19728_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .X(_02147_));
 sky130_fd_sc_hd__nand2_2 _19729_ (.A(net59),
    .B(_10653_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand4_1 _19730_ (.A(_10542_),
    .B(_10639_),
    .C(_10924_),
    .D(_01653_),
    .Y(_02149_));
 sky130_fd_sc_hd__o41ai_4 _19731_ (.A1(net25),
    .A2(\load_store_unit_i.lsu_err_q ),
    .A3(\load_store_unit_i.data_we_q ),
    .A4(_02148_),
    .B1(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__and3_4 _19732_ (.A(net3829),
    .B(net3828),
    .C(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_535 ();
 sky130_fd_sc_hd__nand2_8 _19734_ (.A(_02147_),
    .B(_02151_),
    .Y(_02153_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_533 ();
 sky130_fd_sc_hd__nand2_1 _19737_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .B(_02153_),
    .Y(_02156_));
 sky130_fd_sc_hd__o21ai_0 _19738_ (.A1(_02145_),
    .A2(_02153_),
    .B1(_02156_),
    .Y(_00514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_530 ();
 sky130_fd_sc_hd__mux4_2 _19742_ (.A0(net58),
    .A1(\load_store_unit_i.rdata_q[9] ),
    .A2(\load_store_unit_i.rdata_q[17] ),
    .A3(net38),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(net3822),
    .X(_02160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_529 ();
 sky130_fd_sc_hd__mux2i_1 _19744_ (.A0(net44),
    .A1(net38),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02162_));
 sky130_fd_sc_hd__mux2_1 _19745_ (.A0(net58),
    .A1(net35),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_02163_));
 sky130_fd_sc_hd__nor2_1 _19746_ (.A(net3822),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _19747_ (.A1(net3822),
    .A2(_02162_),
    .B1(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__a22oi_1 _19748_ (.A1(_01670_),
    .A2(_02160_),
    .B1(_02165_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .Y(_02166_));
 sky130_fd_sc_hd__nand3_4 _19749_ (.A(net3472),
    .B(_01669_),
    .C(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_526 ();
 sky130_fd_sc_hd__xnor2_4 _19753_ (.A(_10547_),
    .B(_02012_),
    .Y(_02171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_525 ();
 sky130_fd_sc_hd__mux2i_2 _19755_ (.A0(_02073_),
    .A1(_02066_),
    .S(net3578),
    .Y(_02173_));
 sky130_fd_sc_hd__mux2i_1 _19756_ (.A0(_02086_),
    .A1(_02071_),
    .S(net3578),
    .Y(_02174_));
 sky130_fd_sc_hd__mux2i_1 _19757_ (.A0(_02173_),
    .A1(_02174_),
    .S(net3558),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _19758_ (.A(net3578),
    .B(_02068_),
    .Y(_02176_));
 sky130_fd_sc_hd__a21oi_2 _19759_ (.A1(_02077_),
    .A2(net3578),
    .B1(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _19760_ (.A(_02077_),
    .B(net3558),
    .Y(_02178_));
 sky130_fd_sc_hd__a21o_4 _19761_ (.A1(net3558),
    .A2(_02177_),
    .B1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2i_1 _19762_ (.A0(_02175_),
    .A1(_02179_),
    .S(_02056_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _19763_ (.A(net3557),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_4 _19764_ (.A(net3560),
    .B(_02077_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_2 _19765_ (.A(_02181_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__and2_4 _19766_ (.A(_02124_),
    .B(_02126_),
    .X(_02184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_524 ();
 sky130_fd_sc_hd__nand2_1 _19768_ (.A(net3618),
    .B(net3617),
    .Y(_02186_));
 sky130_fd_sc_hd__xnor2_1 _19769_ (.A(net3726),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_523 ();
 sky130_fd_sc_hd__o221ai_1 _19771_ (.A1(net3618),
    .A2(net3617),
    .B1(_02184_),
    .B2(_02187_),
    .C1(_02137_),
    .Y(_02189_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_520 ();
 sky130_fd_sc_hd__mux2i_1 _19775_ (.A0(_02082_),
    .A1(_02085_),
    .S(net3619),
    .Y(_02193_));
 sky130_fd_sc_hd__mux2i_1 _19776_ (.A0(_02193_),
    .A1(_02043_),
    .S(net3578),
    .Y(_02194_));
 sky130_fd_sc_hd__mux2i_2 _19777_ (.A0(_02088_),
    .A1(_02093_),
    .S(net3619),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2i_1 _19778_ (.A0(_02094_),
    .A1(_02081_),
    .S(net3619),
    .Y(_02196_));
 sky130_fd_sc_hd__mux2i_1 _19779_ (.A0(_02195_),
    .A1(_02196_),
    .S(net3578),
    .Y(_02197_));
 sky130_fd_sc_hd__mux2i_2 _19780_ (.A0(_02194_),
    .A1(_02197_),
    .S(net3558),
    .Y(_02198_));
 sky130_fd_sc_hd__mux2i_2 _19781_ (.A0(_02100_),
    .A1(_02102_),
    .S(net3619),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _19782_ (.A(net3621),
    .B(net3603),
    .Y(_02200_));
 sky130_fd_sc_hd__mux2_8 _19783_ (.A0(_09310_),
    .A1(_09520_),
    .S(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _19784_ (.A0(_02199_),
    .A1(_02201_),
    .S(net3578),
    .X(_02202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_519 ();
 sky130_fd_sc_hd__mux2i_2 _19786_ (.A0(_02110_),
    .A1(_02112_),
    .S(net3619),
    .Y(_02204_));
 sky130_fd_sc_hd__mux2i_2 _19787_ (.A0(_02114_),
    .A1(_02099_),
    .S(net3619),
    .Y(_02205_));
 sky130_fd_sc_hd__mux2i_1 _19788_ (.A0(_02204_),
    .A1(_02205_),
    .S(net3578),
    .Y(_02206_));
 sky130_fd_sc_hd__nand2_1 _19789_ (.A(net3558),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__o21ai_0 _19790_ (.A1(net3558),
    .A2(_02202_),
    .B1(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _19791_ (.A(net3559),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__o21ai_2 _19792_ (.A1(net3559),
    .A2(_02198_),
    .B1(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_518 ();
 sky130_fd_sc_hd__mux2i_1 _19794_ (.A0(_02048_),
    .A1(_02028_),
    .S(net3578),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2b_1 _19795_ (.A_N(net3578),
    .B(_02035_),
    .Y(_02213_));
 sky130_fd_sc_hd__o211ai_1 _19796_ (.A1(net3621),
    .A2(_02058_),
    .B1(net3578),
    .C1(_02055_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_2 _19797_ (.A(_02213_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _19798_ (.A(net3558),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21oi_2 _19799_ (.A1(net3558),
    .A2(_02212_),
    .B1(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _19800_ (.A(net3559),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__o21ai_1 _19801_ (.A1(_02077_),
    .A2(net3559),
    .B1(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__nor2_1 _19802_ (.A(net3560),
    .B(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__a21oi_4 _19803_ (.A1(net3560),
    .A2(_02210_),
    .B1(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _19804_ (.A(net3602),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__o211ai_1 _19805_ (.A1(_02020_),
    .A2(_02183_),
    .B1(_02189_),
    .C1(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__a21oi_2 _19806_ (.A1(net3520),
    .A2(_02006_),
    .B1(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__nor3_4 _19807_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .C(_01999_),
    .Y(_02225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_517 ();
 sky130_fd_sc_hd__nor3_1 _19809_ (.A(_01775_),
    .B(_01871_),
    .C(_01872_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand3_1 _19810_ (.A(_01775_),
    .B(_01761_),
    .C(_01767_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand3_1 _19811_ (.A(_01875_),
    .B(_01869_),
    .C(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__o21ba_4 _19812_ (.A1(_01755_),
    .A2(_02227_),
    .B1_N(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__nor2_1 _19813_ (.A(net3652),
    .B(_01690_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _19814_ (.A(net3654),
    .B(_01745_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor2_2 _19815_ (.A(net3659),
    .B(_01713_),
    .Y(_02233_));
 sky130_fd_sc_hd__xnor2_1 _19816_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_1 _19817_ (.A(_02231_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__o31ai_4 _19818_ (.A1(_09961_),
    .A2(_09982_),
    .A3(net3761),
    .B1(_01842_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand2_1 _19819_ (.A(_01802_),
    .B(net3637),
    .Y(_02237_));
 sky130_fd_sc_hd__mux2_1 _19820_ (.A0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .S(_10740_),
    .X(_02238_));
 sky130_fd_sc_hd__a22oi_2 _19821_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net3759),
    .B1(_02238_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_02239_));
 sky130_fd_sc_hd__mux2_8 _19822_ (.A0(net3705),
    .A1(_10088_),
    .S(_01685_),
    .X(_02240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_516 ();
 sky130_fd_sc_hd__or3_4 _19824_ (.A(_01711_),
    .B(_02239_),
    .C(_02240_),
    .X(_02242_));
 sky130_fd_sc_hd__or2_4 _19825_ (.A(_01743_),
    .B(_01744_),
    .X(_02243_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_515 ();
 sky130_fd_sc_hd__a41o_1 _19827_ (.A1(_01802_),
    .A2(_01794_),
    .A3(_02243_),
    .A4(net3637),
    .B1(_01841_),
    .X(_02245_));
 sky130_fd_sc_hd__o221ai_1 _19828_ (.A1(_01844_),
    .A2(_01845_),
    .B1(_02237_),
    .B2(_02242_),
    .C1(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_514 ();
 sky130_fd_sc_hd__o32ai_1 _19830_ (.A1(_01711_),
    .A2(_02239_),
    .A3(_02240_),
    .B1(net3639),
    .B2(_01700_),
    .Y(_02248_));
 sky130_fd_sc_hd__o21ai_2 _19831_ (.A1(_01711_),
    .A2(_02240_),
    .B1(_02239_),
    .Y(_02249_));
 sky130_fd_sc_hd__mux2i_1 _19832_ (.A0(_02237_),
    .A1(_02248_),
    .S(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_2 _19833_ (.A(_01700_),
    .B(net3639),
    .Y(_02251_));
 sky130_fd_sc_hd__o311ai_0 _19834_ (.A1(_01711_),
    .A2(_02239_),
    .A3(_02240_),
    .B1(net3637),
    .C1(_01802_),
    .Y(_02252_));
 sky130_fd_sc_hd__mux2i_1 _19835_ (.A0(_02251_),
    .A1(_02252_),
    .S(_02249_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _19836_ (.A(_01802_),
    .B(_02243_),
    .Y(_02254_));
 sky130_fd_sc_hd__a21oi_1 _19837_ (.A1(_01794_),
    .A2(net3637),
    .B1(_01841_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand3_1 _19838_ (.A(_01794_),
    .B(_01841_),
    .C(net3637),
    .Y(_02256_));
 sky130_fd_sc_hd__o221ai_1 _19839_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02242_),
    .B2(_02251_),
    .C1(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__o22ai_2 _19840_ (.A1(_02246_),
    .A2(_02250_),
    .B1(_02253_),
    .B2(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__xnor2_2 _19841_ (.A(_02235_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__maj3_4 _19842_ (.A(_01846_),
    .B(_01850_),
    .C(_01854_),
    .X(_02260_));
 sky130_fd_sc_hd__nand2_2 _19843_ (.A(_01815_),
    .B(_01780_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_2 _19844_ (.A(_01689_),
    .B(_01765_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_2 _19845_ (.A(_01693_),
    .B(_01775_),
    .Y(_02263_));
 sky130_fd_sc_hd__xnor3_1 _19846_ (.A(_02261_),
    .B(_02262_),
    .C(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__maj3_1 _19847_ (.A(net3606),
    .B(net3605),
    .C(_01859_),
    .X(_02265_));
 sky130_fd_sc_hd__maj3_1 _19848_ (.A(_01851_),
    .B(_01852_),
    .C(_01853_),
    .X(_02266_));
 sky130_fd_sc_hd__xnor3_1 _19849_ (.A(_02264_),
    .B(_02265_),
    .C(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__xnor2_1 _19850_ (.A(_02260_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__xnor2_1 _19851_ (.A(_02259_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__mux2_8 _19852_ (.A0(net3706),
    .A1(net3684),
    .S(_01681_),
    .X(_02270_));
 sky130_fd_sc_hd__nand2_1 _19853_ (.A(_01771_),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _19854_ (.A(net3648),
    .B(_01867_),
    .Y(_02272_));
 sky130_fd_sc_hd__xnor2_1 _19855_ (.A(_02271_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__maj3_2 _19856_ (.A(_01856_),
    .B(_01860_),
    .C(_01861_),
    .X(_02274_));
 sky130_fd_sc_hd__xnor2_1 _19857_ (.A(_02273_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__maj3_2 _19858_ (.A(_01855_),
    .B(_01862_),
    .C(_01863_),
    .X(_02276_));
 sky130_fd_sc_hd__xor2_1 _19859_ (.A(_02275_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__xnor2_1 _19860_ (.A(_02277_),
    .B(_02269_),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_1 _19861_ (.A(_02230_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2_1 _19862_ (.A(_01865_),
    .B(_01878_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _19863_ (.A(_01865_),
    .B(_01878_),
    .Y(_02281_));
 sky130_fd_sc_hd__a21oi_2 _19864_ (.A1(_01877_),
    .A2(_02280_),
    .B1(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__xnor2_1 _19865_ (.A(_02279_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__o22a_1 _19866_ (.A1(_01838_),
    .A2(_01880_),
    .B1(_01885_),
    .B2(_01925_),
    .X(_02284_));
 sky130_fd_sc_hd__a21oi_1 _19867_ (.A1(_01838_),
    .A2(_01880_),
    .B1(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__xor2_2 _19868_ (.A(net3521),
    .B(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__xnor2_1 _19869_ (.A(_01885_),
    .B(_01925_),
    .Y(_02287_));
 sky130_fd_sc_hd__or3_4 _19870_ (.A(net3523),
    .B(net3531),
    .C(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__xnor2_4 _19871_ (.A(_02286_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _19872_ (.A(_02225_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__a21oi_2 _19873_ (.A1(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .A2(_02225_),
    .B1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_513 ();
 sky130_fd_sc_hd__nand2_1 _19875_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .Y(_02293_));
 sky130_fd_sc_hd__o21ai_4 _19876_ (.A1(net3937),
    .A2(_02291_),
    .B1(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_2 _19877_ (.A(_07857_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__o2111ai_4 _19878_ (.A1(net3755),
    .A2(_02224_),
    .B1(_02295_),
    .C1(_11724_),
    .D1(_01655_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_8 _19879_ (.A(_02167_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_512 ();
 sky130_fd_sc_hd__nand2_1 _19881_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .B(_02153_),
    .Y(_02299_));
 sky130_fd_sc_hd__o21ai_0 _19882_ (.A1(_02153_),
    .A2(_02297_),
    .B1(_02299_),
    .Y(_00515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_511 ();
 sky130_fd_sc_hd__mux4_2 _19884_ (.A0(net28),
    .A1(net36),
    .A2(net45),
    .A3(net49),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux4_2 _19885_ (.A0(net28),
    .A1(\load_store_unit_i.rdata_q[10] ),
    .A2(\load_store_unit_i.rdata_q[18] ),
    .A3(net49),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02302_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_510 ();
 sky130_fd_sc_hd__a22oi_1 _19887_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02301_),
    .B1(_02302_),
    .B2(_01670_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand3_4 _19888_ (.A(net3472),
    .B(_01669_),
    .C(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_509 ();
 sky130_fd_sc_hd__a21o_1 _19890_ (.A1(net3606),
    .A2(net3605),
    .B1(_01859_),
    .X(_02307_));
 sky130_fd_sc_hd__o21ai_4 _19891_ (.A1(net3606),
    .A2(net3605),
    .B1(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__xnor2_1 _19892_ (.A(_02262_),
    .B(_02263_),
    .Y(_02309_));
 sky130_fd_sc_hd__xnor2_1 _19893_ (.A(_02261_),
    .B(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__a21o_1 _19894_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01851_),
    .X(_02311_));
 sky130_fd_sc_hd__o21ai_2 _19895_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__maj3_2 _19896_ (.A(_02259_),
    .B(_02310_),
    .C(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__o2111a_1 _19897_ (.A1(_02260_),
    .A2(_02308_),
    .B1(_02312_),
    .C1(_02310_),
    .D1(_02259_),
    .X(_02314_));
 sky130_fd_sc_hd__a31o_4 _19898_ (.A1(_02260_),
    .A2(_02308_),
    .A3(_02313_),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__a2111o_1 _19899_ (.A1(_02260_),
    .A2(_02308_),
    .B1(_02312_),
    .C1(_02310_),
    .D1(_02259_),
    .X(_02316_));
 sky130_fd_sc_hd__o31ai_1 _19900_ (.A1(_02260_),
    .A2(_02308_),
    .A3(_02313_),
    .B1(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__mux2i_4 _19901_ (.A0(net3706),
    .A1(_10057_),
    .S(_01681_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_2 _19902_ (.A(net3648),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__mux2_8 _19903_ (.A0(net333),
    .A1(_10131_),
    .S(net3760),
    .X(_02320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_508 ();
 sky130_fd_sc_hd__a22oi_1 _19905_ (.A1(_01762_),
    .A2(_02319_),
    .B1(_02320_),
    .B2(_01869_),
    .Y(_02322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_507 ();
 sky130_fd_sc_hd__mux2i_2 _19907_ (.A0(net333),
    .A1(_10131_),
    .S(net3760),
    .Y(_02324_));
 sky130_fd_sc_hd__o22ai_1 _19908_ (.A1(net3648),
    .A2(_02318_),
    .B1(net3635),
    .B2(_01762_),
    .Y(_02325_));
 sky130_fd_sc_hd__nand3_1 _19909_ (.A(net3644),
    .B(_02319_),
    .C(_02320_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_1 _19910_ (.A(_01762_),
    .B(_02319_),
    .Y(_02327_));
 sky130_fd_sc_hd__a211oi_1 _19911_ (.A1(net3644),
    .A2(_02320_),
    .B1(net3638),
    .C1(_01689_),
    .Y(_02328_));
 sky130_fd_sc_hd__a32oi_2 _19912_ (.A1(net3638),
    .A2(_02325_),
    .A3(_02326_),
    .B1(_02327_),
    .B2(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__o21ai_4 _19913_ (.A1(_01886_),
    .A2(_02322_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand2_2 _19914_ (.A(_02249_),
    .B(_02248_),
    .Y(_02331_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .S(_10740_),
    .X(_02332_));
 sky130_fd_sc_hd__a22oi_2 _19916_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net3759),
    .B1(_02332_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_02333_));
 sky130_fd_sc_hd__mux2_8 _19917_ (.A0(net400),
    .A1(_10157_),
    .S(_01685_),
    .X(_02334_));
 sky130_fd_sc_hd__nor2_2 _19918_ (.A(net3651),
    .B(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__nor2_1 _19919_ (.A(_01700_),
    .B(_02240_),
    .Y(_02336_));
 sky130_fd_sc_hd__xor3_1 _19920_ (.A(_02333_),
    .B(_02335_),
    .C(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__nor2_1 _19921_ (.A(net3654),
    .B(_01843_),
    .Y(_02338_));
 sky130_fd_sc_hd__nor2_2 _19922_ (.A(net3659),
    .B(_01745_),
    .Y(_02339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_506 ();
 sky130_fd_sc_hd__nor2_1 _19924_ (.A(net417),
    .B(_01713_),
    .Y(_02341_));
 sky130_fd_sc_hd__xnor3_1 _19925_ (.A(_02338_),
    .B(_02339_),
    .C(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__xnor2_1 _19926_ (.A(_02337_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__xor2_1 _19927_ (.A(_02331_),
    .B(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__nor2_1 _19928_ (.A(net3652),
    .B(net3643),
    .Y(_02345_));
 sky130_fd_sc_hd__nor2_1 _19929_ (.A(_01693_),
    .B(_01759_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _19930_ (.A(net3660),
    .B(_01765_),
    .Y(_02347_));
 sky130_fd_sc_hd__xor2_1 _19931_ (.A(_02346_),
    .B(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__xnor2_1 _19932_ (.A(_02345_),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__maj3_4 _19933_ (.A(_02231_),
    .B(_02232_),
    .C(_02233_),
    .X(_02350_));
 sky130_fd_sc_hd__nor2_1 _19934_ (.A(net3660),
    .B(_01759_),
    .Y(_02351_));
 sky130_fd_sc_hd__maj3_4 _19935_ (.A(_02351_),
    .B(_02262_),
    .C(_02263_),
    .X(_02352_));
 sky130_fd_sc_hd__xor2_1 _19936_ (.A(_02350_),
    .B(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__xnor2_1 _19937_ (.A(_02349_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__o21ai_0 _19938_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02256_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_1 _19939_ (.A(_02249_),
    .B(_02242_),
    .Y(_02356_));
 sky130_fd_sc_hd__xnor2_1 _19940_ (.A(_02251_),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__maj3_4 _19941_ (.A(_02235_),
    .B(_02355_),
    .C(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__xnor3_1 _19942_ (.A(_02344_),
    .B(_02354_),
    .C(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__xor2_1 _19943_ (.A(_02330_),
    .B(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__o21ai_2 _19944_ (.A1(_02315_),
    .A2(_02317_),
    .B1(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__a31oi_1 _19945_ (.A1(_02260_),
    .A2(_02308_),
    .A3(_02313_),
    .B1(_02314_),
    .Y(_02362_));
 sky130_fd_sc_hd__o31a_1 _19946_ (.A1(_02260_),
    .A2(_02308_),
    .A3(_02313_),
    .B1(_02316_),
    .X(_02363_));
 sky130_fd_sc_hd__xnor2_1 _19947_ (.A(_02330_),
    .B(_02359_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand3_2 _19948_ (.A(_02362_),
    .B(_02363_),
    .C(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_2 _19949_ (.A(_02273_),
    .B(_02274_),
    .Y(_02366_));
 sky130_fd_sc_hd__maj3_1 _19950_ (.A(_02275_),
    .B(_02276_),
    .C(_02269_),
    .X(_02367_));
 sky130_fd_sc_hd__nor3_1 _19951_ (.A(_02366_),
    .B(_02276_),
    .C(_02269_),
    .Y(_02368_));
 sky130_fd_sc_hd__a21o_4 _19952_ (.A1(_02366_),
    .A2(_02367_),
    .B1(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__a21o_4 _19953_ (.A1(_02361_),
    .A2(_02365_),
    .B1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__nand3_2 _19954_ (.A(_02361_),
    .B(_02365_),
    .C(_02369_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _19955_ (.A(_02230_),
    .B(net3543),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _19956_ (.A(_02230_),
    .B(net3543),
    .Y(_02373_));
 sky130_fd_sc_hd__o21a_4 _19957_ (.A1(_02372_),
    .A2(_02282_),
    .B1(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__a21oi_1 _19958_ (.A1(_02370_),
    .A2(_02371_),
    .B1(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand3_2 _19959_ (.A(_02370_),
    .B(_02371_),
    .C(_02374_),
    .Y(_02376_));
 sky130_fd_sc_hd__nand2b_4 _19960_ (.A_N(_02375_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__xnor2_1 _19961_ (.A(_01865_),
    .B(_01878_),
    .Y(_02378_));
 sky130_fd_sc_hd__mux2_1 _19962_ (.A0(_02378_),
    .A1(_02280_),
    .S(_01877_),
    .X(_02379_));
 sky130_fd_sc_hd__nand2_1 _19963_ (.A(_01877_),
    .B(_02281_),
    .Y(_02380_));
 sky130_fd_sc_hd__mux2_2 _19964_ (.A0(_02379_),
    .A1(_02380_),
    .S(_02279_),
    .X(_02381_));
 sky130_fd_sc_hd__o32a_1 _19965_ (.A1(_01881_),
    .A2(_01997_),
    .A3(_02283_),
    .B1(_02381_),
    .B2(_01838_),
    .X(_02382_));
 sky130_fd_sc_hd__xor2_4 _19966_ (.A(_02377_),
    .B(net3518),
    .X(_02383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_505 ();
 sky130_fd_sc_hd__mux2i_2 _19968_ (.A0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A1(_02383_),
    .S(_02000_),
    .Y(_02385_));
 sky130_fd_sc_hd__nand2_1 _19969_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .Y(_02386_));
 sky130_fd_sc_hd__o21ai_4 _19970_ (.A1(net3937),
    .A2(_02385_),
    .B1(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand2_1 _19971_ (.A(net151),
    .B(_02006_),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _19972_ (.A(_02177_),
    .Y(_02389_));
 sky130_fd_sc_hd__mux2i_4 _19973_ (.A0(_02389_),
    .A1(_02173_),
    .S(net3558),
    .Y(_02390_));
 sky130_fd_sc_hd__o21ai_2 _19974_ (.A1(_02056_),
    .A2(_02390_),
    .B1(_02078_),
    .Y(_02391_));
 sky130_fd_sc_hd__mux2i_1 _19975_ (.A0(_02106_),
    .A1(_02092_),
    .S(net3578),
    .Y(_02392_));
 sky130_fd_sc_hd__mux2_1 _19976_ (.A0(_02115_),
    .A1(_02101_),
    .S(net3578),
    .X(_02393_));
 sky130_fd_sc_hd__nand2_1 _19977_ (.A(net3558),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__o21ai_0 _19978_ (.A1(net3558),
    .A2(_02392_),
    .B1(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__mux2i_1 _19979_ (.A0(_02095_),
    .A1(_02083_),
    .S(net3578),
    .Y(_02396_));
 sky130_fd_sc_hd__mux2i_1 _19980_ (.A0(_02174_),
    .A1(_02396_),
    .S(net3558),
    .Y(_02397_));
 sky130_fd_sc_hd__nand2b_1 _19981_ (.A_N(_02397_),
    .B(_02056_),
    .Y(_02398_));
 sky130_fd_sc_hd__o211ai_1 _19982_ (.A1(_02056_),
    .A2(_02395_),
    .B1(_02398_),
    .C1(net3560),
    .Y(_02399_));
 sky130_fd_sc_hd__o21ai_2 _19983_ (.A1(net3560),
    .A2(_02391_),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__mux2i_2 _19984_ (.A0(_02212_),
    .A1(_02194_),
    .S(net3558),
    .Y(_02401_));
 sky130_fd_sc_hd__a21oi_1 _19985_ (.A1(net3558),
    .A2(_02215_),
    .B1(_02178_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _19986_ (.A(net3559),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__a21oi_4 _19987_ (.A1(net3559),
    .A2(_02401_),
    .B1(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__a21oi_2 _19988_ (.A1(net3560),
    .A2(_02404_),
    .B1(_02063_),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_1 _19989_ (.A(_10563_),
    .B(net3592),
    .Y(_02406_));
 sky130_fd_sc_hd__xnor2_1 _19990_ (.A(_02129_),
    .B(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__o21ai_0 _19991_ (.A1(_10563_),
    .A2(net3592),
    .B1(_02137_),
    .Y(_02408_));
 sky130_fd_sc_hd__a21oi_1 _19992_ (.A1(_02127_),
    .A2(_02407_),
    .B1(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__a221oi_2 _19993_ (.A1(net3602),
    .A2(_02400_),
    .B1(_02405_),
    .B2(net3603),
    .C1(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand3_1 _19994_ (.A(net3745),
    .B(_02388_),
    .C(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__o21ai_4 _19995_ (.A1(net3745),
    .A2(_02387_),
    .B1(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand3_4 _19996_ (.A(_11143_),
    .B(net3469),
    .C(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__nand2_8 _19997_ (.A(_02305_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_504 ();
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .B(_02153_),
    .Y(_02416_));
 sky130_fd_sc_hd__o21ai_0 _20000_ (.A1(_02153_),
    .A2(_02414_),
    .B1(_02416_),
    .Y(_00516_));
 sky130_fd_sc_hd__nor2_4 _20001_ (.A(\load_store_unit_i.data_type_q[2] ),
    .B(_10666_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_4 _20002_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02418_));
 sky130_fd_sc_hd__clkinv_8 _20003_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02419_));
 sky130_fd_sc_hd__nor2_4 _20004_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_503 ();
 sky130_fd_sc_hd__a22oi_1 _20006_ (.A1(_02419_),
    .A2(net46),
    .B1(net37),
    .B2(_02420_),
    .Y(_02422_));
 sky130_fd_sc_hd__inv_8 _20007_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_4 _20008_ (.A(_02423_),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02424_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_502 ();
 sky130_fd_sc_hd__a221oi_1 _20010_ (.A1(_02423_),
    .A2(\load_store_unit_i.rdata_q[11] ),
    .B1(_02424_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_02426_));
 sky130_fd_sc_hd__a21oi_1 _20011_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02422_),
    .B1(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_500 ();
 sky130_fd_sc_hd__a21oi_1 _20014_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net52),
    .B1(_02427_),
    .Y(_02430_));
 sky130_fd_sc_hd__nor2_1 _20015_ (.A(_02423_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__a221oi_1 _20016_ (.A1(net29),
    .A2(_02418_),
    .B1(_02427_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .C1(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__o21ai_2 _20017_ (.A1(_02417_),
    .A2(_02432_),
    .B1(_01669_),
    .Y(_02433_));
 sky130_fd_sc_hd__mux2i_1 _20018_ (.A0(_02075_),
    .A1(_02087_),
    .S(net3558),
    .Y(_02434_));
 sky130_fd_sc_hd__mux2i_1 _20019_ (.A0(_02077_),
    .A1(_02070_),
    .S(net3558),
    .Y(_02435_));
 sky130_fd_sc_hd__mux2i_1 _20020_ (.A0(_02434_),
    .A1(_02435_),
    .S(_02056_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _20021_ (.A(net3557),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_2 _20022_ (.A(_02182_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_499 ();
 sky130_fd_sc_hd__nand2_1 _20024_ (.A(_09026_),
    .B(_08988_),
    .Y(_02440_));
 sky130_fd_sc_hd__xnor2_1 _20025_ (.A(_02133_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__o221ai_1 _20026_ (.A1(_09026_),
    .A2(_08988_),
    .B1(_02184_),
    .B2(_02441_),
    .C1(_02137_),
    .Y(_02442_));
 sky130_fd_sc_hd__o21ai_0 _20027_ (.A1(_10600_),
    .A2(_02058_),
    .B1(_02055_),
    .Y(_02443_));
 sky130_fd_sc_hd__mux2i_2 _20028_ (.A0(_02443_),
    .A1(_02039_),
    .S(net3558),
    .Y(_02444_));
 sky130_fd_sc_hd__o21ai_2 _20029_ (.A1(_02056_),
    .A2(_02444_),
    .B1(_02078_),
    .Y(_02445_));
 sky130_fd_sc_hd__mux2i_1 _20030_ (.A0(_02196_),
    .A1(_02193_),
    .S(net3578),
    .Y(_02446_));
 sky130_fd_sc_hd__mux2i_1 _20031_ (.A0(_02049_),
    .A1(_02446_),
    .S(net3558),
    .Y(_02447_));
 sky130_fd_sc_hd__mux2i_1 _20032_ (.A0(_02201_),
    .A1(_02195_),
    .S(net3578),
    .Y(_02448_));
 sky130_fd_sc_hd__mux2i_1 _20033_ (.A0(_02205_),
    .A1(_02199_),
    .S(net3578),
    .Y(_02449_));
 sky130_fd_sc_hd__mux2_1 _20034_ (.A0(_02448_),
    .A1(_02449_),
    .S(net3558),
    .X(_02450_));
 sky130_fd_sc_hd__nand2_1 _20035_ (.A(net3559),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__o211ai_1 _20036_ (.A1(net3559),
    .A2(_02447_),
    .B1(_02451_),
    .C1(net3560),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_2 _20037_ (.A1(net3560),
    .A2(_02445_),
    .B1(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _20038_ (.A(net3602),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__o211ai_1 _20039_ (.A1(_02020_),
    .A2(_02438_),
    .B1(_02442_),
    .C1(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_498 ();
 sky130_fd_sc_hd__a211oi_1 _20041_ (.A1(net152),
    .A2(_02006_),
    .B1(_02455_),
    .C1(net3755),
    .Y(_02457_));
 sky130_fd_sc_hd__a21oi_1 _20042_ (.A1(_02362_),
    .A2(_02363_),
    .B1(_02364_),
    .Y(_02458_));
 sky130_fd_sc_hd__nor3_1 _20043_ (.A(_02315_),
    .B(_02317_),
    .C(_02360_),
    .Y(_02459_));
 sky130_fd_sc_hd__o31a_1 _20044_ (.A1(_02366_),
    .A2(_02458_),
    .A3(_02459_),
    .B1(_02367_),
    .X(_02460_));
 sky130_fd_sc_hd__a21boi_2 _20045_ (.A1(_02361_),
    .A2(_02365_),
    .B1_N(_02366_),
    .Y(_02461_));
 sky130_fd_sc_hd__nand2b_4 _20046_ (.A_N(_02359_),
    .B(_02330_),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_1 _20047_ (.A(_02363_),
    .B(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2b_1 _20048_ (.A(_02330_),
    .B_N(_02359_),
    .Y(_02464_));
 sky130_fd_sc_hd__a22o_4 _20049_ (.A1(_02315_),
    .A2(_02462_),
    .B1(_02464_),
    .B2(_02363_),
    .X(_02465_));
 sky130_fd_sc_hd__o21ai_0 _20050_ (.A1(_01700_),
    .A2(_02240_),
    .B1(_02333_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor3_1 _20051_ (.A(_01700_),
    .B(_02240_),
    .C(_02333_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21oi_1 _20052_ (.A1(_02335_),
    .A2(_02466_),
    .B1(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__nor2_1 _20053_ (.A(net449),
    .B(_02240_),
    .Y(_02469_));
 sky130_fd_sc_hd__nor2_2 _20054_ (.A(_01690_),
    .B(_01745_),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_2 _20055_ (.A(net3659),
    .B(_01843_),
    .Y(_02471_));
 sky130_fd_sc_hd__xnor3_1 _20056_ (.A(_02469_),
    .B(_02470_),
    .C(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__nor2_1 _20057_ (.A(_10204_),
    .B(_01999_),
    .Y(_02473_));
 sky130_fd_sc_hd__a21oi_2 _20058_ (.A1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .A2(_01999_),
    .B1(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__o22ai_4 _20059_ (.A1(_10204_),
    .A2(net3757),
    .B1(_02474_),
    .B2(_01738_),
    .Y(_02475_));
 sky130_fd_sc_hd__mux2_8 _20060_ (.A0(net3702),
    .A1(_10199_),
    .S(_01685_),
    .X(_02476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_497 ();
 sky130_fd_sc_hd__nor2_2 _20062_ (.A(net3651),
    .B(_02476_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_2 _20063_ (.A(_01700_),
    .B(_02334_),
    .Y(_02479_));
 sky130_fd_sc_hd__xor3_1 _20064_ (.A(_02475_),
    .B(_02478_),
    .C(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__xnor3_1 _20065_ (.A(_02468_),
    .B(_02472_),
    .C(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__maj3_1 _20066_ (.A(_02331_),
    .B(_02337_),
    .C(_02342_),
    .X(_02482_));
 sky130_fd_sc_hd__nor4_1 _20067_ (.A(net3652),
    .B(_01693_),
    .C(net3642),
    .D(_01759_),
    .Y(_02483_));
 sky130_fd_sc_hd__o22ai_1 _20068_ (.A1(net3652),
    .A2(net3642),
    .B1(_01759_),
    .B2(_01693_),
    .Y(_02484_));
 sky130_fd_sc_hd__o21ai_1 _20069_ (.A1(_02347_),
    .A2(_02483_),
    .B1(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor4_1 _20070_ (.A(net417),
    .B(net3654),
    .C(_01713_),
    .D(_01843_),
    .Y(_02486_));
 sky130_fd_sc_hd__o22ai_1 _20071_ (.A1(net417),
    .A2(_01713_),
    .B1(_01843_),
    .B2(net3654),
    .Y(_02487_));
 sky130_fd_sc_hd__o21ai_2 _20072_ (.A1(_02339_),
    .A2(_02486_),
    .B1(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _20073_ (.A(net3652),
    .B(_01759_),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _20074_ (.A(net444),
    .B(net3642),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_1 _20075_ (.A(_01693_),
    .B(_01765_),
    .Y(_02491_));
 sky130_fd_sc_hd__xnor3_1 _20076_ (.A(_02489_),
    .B(_02490_),
    .C(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__xor3_1 _20077_ (.A(_02485_),
    .B(_02488_),
    .C(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__xnor2_1 _20078_ (.A(_02482_),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__xor2_1 _20079_ (.A(_02481_),
    .B(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__nor2_1 _20080_ (.A(_02350_),
    .B(_02352_),
    .Y(_02496_));
 sky130_fd_sc_hd__nand2_1 _20081_ (.A(_02350_),
    .B(_02352_),
    .Y(_02497_));
 sky130_fd_sc_hd__o21a_1 _20082_ (.A1(_02349_),
    .A2(_02496_),
    .B1(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__nor2_1 _20083_ (.A(net3648),
    .B(net3635),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _20084_ (.A(net397),
    .B(_01867_),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _20085_ (.A(_01689_),
    .B(_02318_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor3_1 _20086_ (.A(_02499_),
    .B(_02500_),
    .C(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_8 _20087_ (.A0(_08917_),
    .A1(_10010_),
    .S(net3760),
    .X(_02503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_496 ();
 sky130_fd_sc_hd__mux2_8 _20089_ (.A0(_09030_),
    .A1(_10229_),
    .S(_01681_),
    .X(_02505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_495 ();
 sky130_fd_sc_hd__o31ai_1 _20091_ (.A1(net3648),
    .A2(_02318_),
    .A3(net3635),
    .B1(_02505_),
    .Y(_02507_));
 sky130_fd_sc_hd__a32oi_1 _20092_ (.A1(_01886_),
    .A2(_02503_),
    .A3(_02325_),
    .B1(_02507_),
    .B2(net3644),
    .Y(_02508_));
 sky130_fd_sc_hd__o32ai_1 _20093_ (.A1(net3648),
    .A2(_02318_),
    .A3(net3635),
    .B1(net3638),
    .B2(_01689_),
    .Y(_02509_));
 sky130_fd_sc_hd__nor2_1 _20094_ (.A(_01762_),
    .B(_02505_),
    .Y(_02510_));
 sky130_fd_sc_hd__o211ai_1 _20095_ (.A1(_02319_),
    .A2(_02320_),
    .B1(_02509_),
    .C1(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2b_1 _20096_ (.A_N(_02508_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__xnor2_1 _20097_ (.A(_02502_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__nor2_2 _20098_ (.A(_01689_),
    .B(_02324_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _20099_ (.A(_01886_),
    .B(_02320_),
    .Y(_02515_));
 sky130_fd_sc_hd__o211a_1 _20100_ (.A1(_02514_),
    .A2(_02515_),
    .B1(_01869_),
    .C1(_02319_),
    .X(_02516_));
 sky130_fd_sc_hd__inv_1 _20101_ (.A(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__xnor3_1 _20102_ (.A(_02498_),
    .B(_02513_),
    .C(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__maj3_1 _20103_ (.A(_02344_),
    .B(_02354_),
    .C(_02358_),
    .X(_02519_));
 sky130_fd_sc_hd__xor3_1 _20104_ (.A(_02495_),
    .B(_02518_),
    .C(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__o21bai_1 _20105_ (.A1(_02463_),
    .A2(_02465_),
    .B1_N(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__a22oi_1 _20106_ (.A1(_02315_),
    .A2(_02462_),
    .B1(_02464_),
    .B2(_02363_),
    .Y(_02522_));
 sky130_fd_sc_hd__nand3b_1 _20107_ (.A_N(_02463_),
    .B(_02522_),
    .C(_02520_),
    .Y(_02523_));
 sky130_fd_sc_hd__a2bb2oi_2 _20108_ (.A1_N(_02460_),
    .A2_N(_02461_),
    .B1(_02521_),
    .B2(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__and4bb_4 _20109_ (.A_N(_02460_),
    .B_N(_02461_),
    .C(_02521_),
    .D(_02523_),
    .X(_02525_));
 sky130_fd_sc_hd__nor2_2 _20110_ (.A(_02524_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__and2_0 _20111_ (.A(_02370_),
    .B(_02371_),
    .X(_02527_));
 sky130_fd_sc_hd__maj3_1 _20112_ (.A(_02527_),
    .B(_02374_),
    .C(_02382_),
    .X(_02528_));
 sky130_fd_sc_hd__xor2_4 _20113_ (.A(_02526_),
    .B(net3510),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_02000_),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__o21ai_4 _20115_ (.A1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .A2(_02000_),
    .B1(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _20116_ (.A(net3937),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__a211oi_4 _20117_ (.A1(net3937),
    .A2(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B1(net3737),
    .C1(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__o211ai_1 _20118_ (.A1(_02457_),
    .A2(_02533_),
    .B1(_11175_),
    .C1(_01655_),
    .Y(_02534_));
 sky130_fd_sc_hd__o21ai_4 _20119_ (.A1(net3469),
    .A2(_02433_),
    .B1(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_494 ();
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .B(_02153_),
    .Y(_02537_));
 sky130_fd_sc_hd__o21ai_0 _20122_ (.A1(_02153_),
    .A2(net3460),
    .B1(_02537_),
    .Y(_00517_));
 sky130_fd_sc_hd__a22oi_1 _20123_ (.A1(_02419_),
    .A2(net47),
    .B1(net39),
    .B2(_02420_),
    .Y(_02538_));
 sky130_fd_sc_hd__a221oi_1 _20124_ (.A1(_02423_),
    .A2(\load_store_unit_i.rdata_q[12] ),
    .B1(_02424_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_02539_));
 sky130_fd_sc_hd__a21oi_1 _20125_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02538_),
    .B1(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21oi_1 _20126_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net53),
    .B1(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _20127_ (.A(_02423_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__a221oi_1 _20128_ (.A1(net30),
    .A2(_02418_),
    .B1(_02540_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .C1(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21ai_2 _20129_ (.A1(_02417_),
    .A2(_02543_),
    .B1(_01669_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _20130_ (.A(_01838_),
    .B(_02381_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor3_1 _20131_ (.A(net3523),
    .B(net3522),
    .C(net3521),
    .Y(_02546_));
 sky130_fd_sc_hd__a211oi_2 _20132_ (.A1(_02376_),
    .A2(_02545_),
    .B1(_02546_),
    .C1(_02375_),
    .Y(_02547_));
 sky130_fd_sc_hd__or2_0 _20133_ (.A(_01838_),
    .B(_02381_),
    .X(_02548_));
 sky130_fd_sc_hd__a311o_1 _20134_ (.A1(_02527_),
    .A2(_02374_),
    .A3(_02548_),
    .B1(_02524_),
    .C1(_02525_),
    .X(_02549_));
 sky130_fd_sc_hd__or2_4 _20135_ (.A(_02547_),
    .B(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__maj3_1 _20136_ (.A(_02495_),
    .B(_02518_),
    .C(_02519_),
    .X(_02551_));
 sky130_fd_sc_hd__maj3_1 _20137_ (.A(_02499_),
    .B(_02500_),
    .C(_02501_),
    .X(_02552_));
 sky130_fd_sc_hd__nor2_1 _20138_ (.A(_01693_),
    .B(_01867_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _20139_ (.A(net397),
    .B(_02318_),
    .Y(_02554_));
 sky130_fd_sc_hd__xor3_1 _20140_ (.A(_02514_),
    .B(_02553_),
    .C(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__mux2i_4 _20141_ (.A0(_09243_),
    .A1(_10294_),
    .S(net3760),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _20142_ (.A(_01771_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__nor2_1 _20143_ (.A(net3648),
    .B(_02505_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_1 _20144_ (.A(_02557_),
    .B(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__xnor3_1 _20145_ (.A(_02552_),
    .B(_02555_),
    .C(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__a21o_4 _20146_ (.A1(_02502_),
    .A2(_02511_),
    .B1(_02508_),
    .X(_02561_));
 sky130_fd_sc_hd__maj3_2 _20147_ (.A(_02485_),
    .B(_02488_),
    .C(_02492_),
    .X(_02562_));
 sky130_fd_sc_hd__xor3_1 _20148_ (.A(_02560_),
    .B(_02561_),
    .C(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__maj3_4 _20149_ (.A(_02481_),
    .B(_02482_),
    .C(_02493_),
    .X(_02564_));
 sky130_fd_sc_hd__o22ai_1 _20150_ (.A1(net444),
    .A2(net3642),
    .B1(_01765_),
    .B2(_01693_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor4_1 _20151_ (.A(_01693_),
    .B(net444),
    .C(net3642),
    .D(_01765_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _20152_ (.A1(_02489_),
    .A2(_02565_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_2 _20153_ (.A(_01713_),
    .B(_01759_),
    .Y(_02568_));
 sky130_fd_sc_hd__o221ai_1 _20154_ (.A1(net3685),
    .A2(_01708_),
    .B1(_01703_),
    .B2(_01704_),
    .C1(_01764_),
    .Y(_02569_));
 sky130_fd_sc_hd__o221ai_1 _20155_ (.A1(_09704_),
    .A2(_01708_),
    .B1(_01743_),
    .B2(_01744_),
    .C1(_01756_),
    .Y(_02570_));
 sky130_fd_sc_hd__xnor2_2 _20156_ (.A(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__xor2_1 _20157_ (.A(_02568_),
    .B(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__nor4_1 _20158_ (.A(net417),
    .B(net449),
    .C(_01745_),
    .D(_02240_),
    .Y(_02573_));
 sky130_fd_sc_hd__o22ai_1 _20159_ (.A1(net417),
    .A2(_01745_),
    .B1(_02240_),
    .B2(net449),
    .Y(_02574_));
 sky130_fd_sc_hd__o21a_4 _20160_ (.A1(_02471_),
    .A2(_02573_),
    .B1(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__xnor3_1 _20161_ (.A(_02567_),
    .B(_02572_),
    .C(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__maj3_2 _20162_ (.A(_02475_),
    .B(_02478_),
    .C(_02479_),
    .X(_02577_));
 sky130_fd_sc_hd__nor2_1 _20163_ (.A(net449),
    .B(_02334_),
    .Y(_02578_));
 sky130_fd_sc_hd__nor2_1 _20164_ (.A(_01690_),
    .B(_01843_),
    .Y(_02579_));
 sky130_fd_sc_hd__nor2_1 _20165_ (.A(net3659),
    .B(_02240_),
    .Y(_02580_));
 sky130_fd_sc_hd__xor3_1 _20166_ (.A(_02578_),
    .B(_02579_),
    .C(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__o41a_1 _20167_ (.A1(_09196_),
    .A2(_09201_),
    .A3(_09205_),
    .A4(_09210_),
    .B1(net3761),
    .X(_02582_));
 sky130_fd_sc_hd__a21o_4 _20168_ (.A1(net3677),
    .A2(_01685_),
    .B1(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__nor2_1 _20169_ (.A(_01711_),
    .B(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__mux2i_1 _20170_ (.A0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .S(_10740_),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _20171_ (.A(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B(net3759),
    .Y(_02586_));
 sky130_fd_sc_hd__o21ai_4 _20172_ (.A1(_01738_),
    .A2(_02585_),
    .B1(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__nor2_1 _20173_ (.A(_01700_),
    .B(_02476_),
    .Y(_02588_));
 sky130_fd_sc_hd__xor3_1 _20174_ (.A(_02584_),
    .B(_02587_),
    .C(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__xor3_1 _20175_ (.A(_02577_),
    .B(_02581_),
    .C(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__xnor3_1 _20176_ (.A(_02475_),
    .B(_02478_),
    .C(_02479_),
    .X(_02591_));
 sky130_fd_sc_hd__maj3_2 _20177_ (.A(_02468_),
    .B(_02472_),
    .C(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__xnor3_1 _20178_ (.A(_02576_),
    .B(_02590_),
    .C(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__xor3_1 _20179_ (.A(_02563_),
    .B(_02564_),
    .C(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__maj3_2 _20180_ (.A(_02498_),
    .B(_02513_),
    .C(_02517_),
    .X(_02595_));
 sky130_fd_sc_hd__xor2_1 _20181_ (.A(_02594_),
    .B(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__xnor2_1 _20182_ (.A(_02551_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__o21bai_1 _20183_ (.A1(_02363_),
    .A2(_02462_),
    .B1_N(_02520_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _20184_ (.A(_02522_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__nand2_2 _20185_ (.A(_02597_),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__inv_1 _20186_ (.A(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__nor3b_4 _20187_ (.A(_02465_),
    .B(_02597_),
    .C_N(_02598_),
    .Y(_02602_));
 sky130_fd_sc_hd__nor2_2 _20188_ (.A(_02601_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__xnor2_1 _20189_ (.A(_02525_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__xor2_4 _20190_ (.A(_02550_),
    .B(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2i_4 _20191_ (.A0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A1(_02605_),
    .S(_02000_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand2_1 _20192_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .Y(_02607_));
 sky130_fd_sc_hd__o21ai_4 _20193_ (.A1(net3937),
    .A2(_02606_),
    .B1(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__mux2_1 _20194_ (.A0(_02096_),
    .A1(_02107_),
    .S(net3558),
    .X(_02609_));
 sky130_fd_sc_hd__nor2_1 _20195_ (.A(_02016_),
    .B(_02434_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21oi_1 _20196_ (.A1(_02016_),
    .A2(_02609_),
    .B1(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand3_4 _20197_ (.A(_02171_),
    .B(_02055_),
    .C(_02058_),
    .Y(_02612_));
 sky130_fd_sc_hd__nand3_1 _20198_ (.A(_02171_),
    .B(_02016_),
    .C(_02435_),
    .Y(_02613_));
 sky130_fd_sc_hd__o21ai_0 _20199_ (.A1(_02016_),
    .A2(_02612_),
    .B1(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a21oi_2 _20200_ (.A1(net3560),
    .A2(_02611_),
    .B1(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__mux2i_2 _20201_ (.A0(_02444_),
    .A1(_02447_),
    .S(net3559),
    .Y(_02616_));
 sky130_fd_sc_hd__o21ai_2 _20202_ (.A1(net3557),
    .A2(_02616_),
    .B1(_02612_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand2_1 _20203_ (.A(_09214_),
    .B(_09245_),
    .Y(_02618_));
 sky130_fd_sc_hd__xor2_1 _20204_ (.A(_02133_),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__o21ai_0 _20205_ (.A1(_09214_),
    .A2(_09245_),
    .B1(_02137_),
    .Y(_02620_));
 sky130_fd_sc_hd__a21oi_1 _20206_ (.A1(_02127_),
    .A2(_02619_),
    .B1(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__a21oi_1 _20207_ (.A1(net3603),
    .A2(_02617_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21ai_0 _20208_ (.A1(_02057_),
    .A2(_02615_),
    .B1(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21oi_1 _20209_ (.A1(net3514),
    .A2(_02006_),
    .B1(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__nand2_2 _20210_ (.A(net3745),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__o21ai_4 _20211_ (.A1(net3745),
    .A2(_02608_),
    .B1(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand3_4 _20212_ (.A(_11195_),
    .B(_01655_),
    .C(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__o21ai_4 _20213_ (.A1(net3469),
    .A2(_02544_),
    .B1(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_493 ();
 sky130_fd_sc_hd__nand2_1 _20215_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .B(_02153_),
    .Y(_02630_));
 sky130_fd_sc_hd__o21ai_0 _20216_ (.A1(_02153_),
    .A2(_02628_),
    .B1(_02630_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand3_1 _20217_ (.A(net3822),
    .B(_02419_),
    .C(net48),
    .Y(_02631_));
 sky130_fd_sc_hd__nand3_1 _20218_ (.A(_02423_),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .C(net40),
    .Y(_02632_));
 sky130_fd_sc_hd__a221oi_1 _20219_ (.A1(_02423_),
    .A2(\load_store_unit_i.rdata_q[13] ),
    .B1(_02424_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_02633_));
 sky130_fd_sc_hd__a31oi_1 _20220_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02631_),
    .A3(_02632_),
    .B1(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_492 ();
 sky130_fd_sc_hd__a21oi_1 _20222_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net54),
    .B1(_02634_),
    .Y(_02636_));
 sky130_fd_sc_hd__nor2_1 _20223_ (.A(_02423_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__a221oi_1 _20224_ (.A1(net31),
    .A2(_02418_),
    .B1(_02634_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .C1(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__o21ai_0 _20225_ (.A1(_02417_),
    .A2(_02638_),
    .B1(_01669_),
    .Y(_02639_));
 sky130_fd_sc_hd__o21bai_2 _20226_ (.A1(_02524_),
    .A2(_02528_),
    .B1_N(_02525_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_4 _20227_ (.A(_02603_),
    .B(net3499),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_1 _20228_ (.A(_02594_),
    .B(_02595_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor2_1 _20229_ (.A(_02594_),
    .B(_02595_),
    .Y(_02643_));
 sky130_fd_sc_hd__a21o_4 _20230_ (.A1(_02551_),
    .A2(_02642_),
    .B1(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__nor2_1 _20231_ (.A(_01705_),
    .B(_01765_),
    .Y(_02645_));
 sky130_fd_sc_hd__nor2_1 _20232_ (.A(_01775_),
    .B(_01745_),
    .Y(_02646_));
 sky130_fd_sc_hd__maj3_1 _20233_ (.A(_02645_),
    .B(_02568_),
    .C(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__nand2_1 _20234_ (.A(_01757_),
    .B(_02236_),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_1 _20235_ (.A(_01780_),
    .B(_02243_),
    .Y(_02649_));
 sky130_fd_sc_hd__nand2b_2 _20236_ (.A_N(_01713_),
    .B(_01783_),
    .Y(_02650_));
 sky130_fd_sc_hd__xnor3_1 _20237_ (.A(_02648_),
    .B(_02649_),
    .C(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__maj3_1 _20238_ (.A(_02578_),
    .B(_02579_),
    .C(_02580_),
    .X(_02652_));
 sky130_fd_sc_hd__xor3_1 _20239_ (.A(_02647_),
    .B(_02651_),
    .C(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__maj3_1 _20240_ (.A(_02584_),
    .B(_02587_),
    .C(_02588_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_8 _20241_ (.A0(net3698),
    .A1(_10332_),
    .S(net3758),
    .X(_02655_));
 sky130_fd_sc_hd__or2_4 _20242_ (.A(_01711_),
    .B(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__a2111oi_2 _20243_ (.A1(net3677),
    .A2(_01685_),
    .B1(_02582_),
    .C1(_01698_),
    .D1(net443),
    .Y(_02657_));
 sky130_fd_sc_hd__mux2i_1 _20244_ (.A0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .S(_10740_),
    .Y(_02658_));
 sky130_fd_sc_hd__nand2_1 _20245_ (.A(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .B(net3759),
    .Y(_02659_));
 sky130_fd_sc_hd__o21ai_4 _20246_ (.A1(_01738_),
    .A2(_02658_),
    .B1(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__xor2_1 _20247_ (.A(_02657_),
    .B(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__xor2_1 _20248_ (.A(_02656_),
    .B(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__nor2_1 _20249_ (.A(net3654),
    .B(_02476_),
    .Y(_02663_));
 sky130_fd_sc_hd__nor2_1 _20250_ (.A(_01690_),
    .B(_02240_),
    .Y(_02664_));
 sky130_fd_sc_hd__nor2_1 _20251_ (.A(net3659),
    .B(_02334_),
    .Y(_02665_));
 sky130_fd_sc_hd__xnor3_1 _20252_ (.A(_02663_),
    .B(_02664_),
    .C(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__xor3_1 _20253_ (.A(_02654_),
    .B(_02662_),
    .C(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__maj3_1 _20254_ (.A(_02577_),
    .B(_02581_),
    .C(_02589_),
    .X(_02668_));
 sky130_fd_sc_hd__xor3_1 _20255_ (.A(_02653_),
    .B(_02667_),
    .C(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__o21ai_0 _20256_ (.A1(_02471_),
    .A2(_02573_),
    .B1(_02574_),
    .Y(_02670_));
 sky130_fd_sc_hd__maj3_1 _20257_ (.A(_02567_),
    .B(_02572_),
    .C(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__maj3_2 _20258_ (.A(_02514_),
    .B(_02553_),
    .C(_02554_),
    .X(_02672_));
 sky130_fd_sc_hd__o21ai_2 _20259_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_02503_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_01815_),
    .B(_02320_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand2_1 _20261_ (.A(_01818_),
    .B(_02270_),
    .Y(_02675_));
 sky130_fd_sc_hd__xnor3_1 _20262_ (.A(_02673_),
    .B(_02674_),
    .C(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_2 _20263_ (.A(_01778_),
    .B(_02556_),
    .Y(_02677_));
 sky130_fd_sc_hd__nor2_1 _20264_ (.A(net3657),
    .B(_02505_),
    .Y(_02678_));
 sky130_fd_sc_hd__nor3b_4 _20265_ (.A(_10345_),
    .B(_10353_),
    .C_N(_10359_),
    .Y(_02679_));
 sky130_fd_sc_hd__mux2_8 _20266_ (.A0(_09149_),
    .A1(_02679_),
    .S(net3760),
    .X(_02680_));
 sky130_fd_sc_hd__nor2_1 _20267_ (.A(_01762_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor3_1 _20268_ (.A(_02677_),
    .B(_02678_),
    .C(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__xnor3_1 _20269_ (.A(_02672_),
    .B(_02676_),
    .C(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__maj3_4 _20270_ (.A(_02552_),
    .B(_02555_),
    .C(_02559_),
    .X(_02684_));
 sky130_fd_sc_hd__xnor3_1 _20271_ (.A(_02671_),
    .B(_02683_),
    .C(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__xnor3_1 _20272_ (.A(_02577_),
    .B(_02581_),
    .C(_02589_),
    .X(_02686_));
 sky130_fd_sc_hd__maj3_4 _20273_ (.A(_02576_),
    .B(_02686_),
    .C(_02592_),
    .X(_02687_));
 sky130_fd_sc_hd__xnor3_1 _20274_ (.A(_02669_),
    .B(_02685_),
    .C(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__maj3_4 _20275_ (.A(_02563_),
    .B(_02564_),
    .C(_02593_),
    .X(_02689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_491 ();
 sky130_fd_sc_hd__nor3_4 _20277_ (.A(_01762_),
    .B(_02505_),
    .C(_02677_),
    .Y(_02691_));
 sky130_fd_sc_hd__maj3_4 _20278_ (.A(_02560_),
    .B(_02561_),
    .C(_02562_),
    .X(_02692_));
 sky130_fd_sc_hd__xnor2_1 _20279_ (.A(_02691_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__xnor2_1 _20280_ (.A(_02689_),
    .B(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__xnor2_1 _20281_ (.A(_02688_),
    .B(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__xor2_2 _20282_ (.A(_02644_),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__xnor2_2 _20283_ (.A(_02602_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__xor2_4 _20284_ (.A(_02641_),
    .B(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__mux2i_4 _20285_ (.A0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .A1(_02698_),
    .S(_02000_),
    .Y(_02699_));
 sky130_fd_sc_hd__nand2_1 _20286_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .Y(_02700_));
 sky130_fd_sc_hd__o21ai_4 _20287_ (.A1(net3937),
    .A2(_02699_),
    .B1(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__nand2_8 _20288_ (.A(net336),
    .B(_10937_),
    .Y(_02702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_490 ();
 sky130_fd_sc_hd__nand2_1 _20290_ (.A(net3558),
    .B(_02202_),
    .Y(_02704_));
 sky130_fd_sc_hd__o21ai_1 _20291_ (.A1(net3558),
    .A2(_02197_),
    .B1(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_1 _20292_ (.A(net3559),
    .B(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand2_1 _20293_ (.A(_02056_),
    .B(_02401_),
    .Y(_02707_));
 sky130_fd_sc_hd__nand2_1 _20294_ (.A(_02706_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__a21oi_1 _20295_ (.A1(net3559),
    .A2(net3558),
    .B1(_02077_),
    .Y(_02709_));
 sky130_fd_sc_hd__a31oi_4 _20296_ (.A1(net3559),
    .A2(net3558),
    .A3(_02215_),
    .B1(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_1 _20297_ (.A(net3560),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a21oi_2 _20298_ (.A1(net3560),
    .A2(_02708_),
    .B1(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_1 _20299_ (.A(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__mux2i_2 _20300_ (.A0(_02390_),
    .A1(_02397_),
    .S(_02016_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21ai_1 _20301_ (.A1(net3557),
    .A2(_02714_),
    .B1(_02612_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2_1 _20302_ (.A(_09158_),
    .B(net3591),
    .Y(_02716_));
 sky130_fd_sc_hd__xor2_1 _20303_ (.A(_02133_),
    .B(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__o21ai_0 _20304_ (.A1(_09158_),
    .A2(net3591),
    .B1(_02137_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21oi_1 _20305_ (.A1(_02127_),
    .A2(_02717_),
    .B1(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__a221oi_1 _20306_ (.A1(net3602),
    .A2(_02713_),
    .B1(_02715_),
    .B2(net3603),
    .C1(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__o211ai_1 _20307_ (.A1(net3498),
    .A2(_02702_),
    .B1(_02720_),
    .C1(net3745),
    .Y(_02721_));
 sky130_fd_sc_hd__o21ai_4 _20308_ (.A1(net3745),
    .A2(_02701_),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__nand3_4 _20309_ (.A(_11212_),
    .B(_01655_),
    .C(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__o21ai_2 _20310_ (.A1(net3469),
    .A2(_02639_),
    .B1(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__nand2_1 _20312_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .B(_02153_),
    .Y(_02726_));
 sky130_fd_sc_hd__o21ai_0 _20313_ (.A1(_02153_),
    .A2(net3453),
    .B1(_02726_),
    .Y(_00519_));
 sky130_fd_sc_hd__mux4_2 _20314_ (.A0(net32),
    .A1(net41),
    .A2(net50),
    .A3(net55),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02727_));
 sky130_fd_sc_hd__mux4_2 _20315_ (.A0(net32),
    .A1(\load_store_unit_i.rdata_q[14] ),
    .A2(\load_store_unit_i.rdata_q[22] ),
    .A3(net55),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02728_));
 sky130_fd_sc_hd__a22oi_1 _20316_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02727_),
    .B1(_02728_),
    .B2(_01670_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand3_2 _20317_ (.A(net3472),
    .B(_01669_),
    .C(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand2_1 _20318_ (.A(_02662_),
    .B(_02666_),
    .Y(_02731_));
 sky130_fd_sc_hd__nor2_1 _20319_ (.A(_02662_),
    .B(_02666_),
    .Y(_02732_));
 sky130_fd_sc_hd__a21o_1 _20320_ (.A1(_02654_),
    .A2(_02731_),
    .B1(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2_1 _20321_ (.A(_02657_),
    .B(_02660_),
    .Y(_02734_));
 sky130_fd_sc_hd__nor2_1 _20322_ (.A(_02657_),
    .B(_02660_),
    .Y(_02735_));
 sky130_fd_sc_hd__a21o_1 _20323_ (.A1(_02656_),
    .A2(_02734_),
    .B1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__nor2_1 _20324_ (.A(net3654),
    .B(_02583_),
    .Y(_02737_));
 sky130_fd_sc_hd__nor2_1 _20325_ (.A(net417),
    .B(_02334_),
    .Y(_02738_));
 sky130_fd_sc_hd__nor2_1 _20326_ (.A(net3658),
    .B(_02476_),
    .Y(_02739_));
 sky130_fd_sc_hd__xnor3_1 _20327_ (.A(_02737_),
    .B(_02738_),
    .C(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2i_1 _20328_ (.A0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .S(_10740_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _20329_ (.A(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B(net3759),
    .Y(_02742_));
 sky130_fd_sc_hd__o21ai_4 _20330_ (.A1(_01738_),
    .A2(_02741_),
    .B1(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__mux2_8 _20331_ (.A0(net3695),
    .A1(_10448_),
    .S(net3758),
    .X(_02744_));
 sky130_fd_sc_hd__nor2_1 _20332_ (.A(_01711_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__nor2_1 _20333_ (.A(_01700_),
    .B(_02655_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor3_1 _20334_ (.A(_02743_),
    .B(_02745_),
    .C(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__xnor3_1 _20335_ (.A(_02736_),
    .B(_02740_),
    .C(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__nor2_1 _20336_ (.A(net3643),
    .B(_02240_),
    .Y(_02749_));
 sky130_fd_sc_hd__nor2_1 _20337_ (.A(_01759_),
    .B(net3639),
    .Y(_02750_));
 sky130_fd_sc_hd__nor2_1 _20338_ (.A(_01745_),
    .B(net3646),
    .Y(_02751_));
 sky130_fd_sc_hd__xnor3_1 _20339_ (.A(_02749_),
    .B(_02750_),
    .C(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__maj3_1 _20340_ (.A(_02648_),
    .B(_02649_),
    .C(_02650_),
    .X(_02753_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__nor4_1 _20343_ (.A(net417),
    .B(net3654),
    .C(_02240_),
    .D(_02476_),
    .Y(_02756_));
 sky130_fd_sc_hd__o22ai_1 _20344_ (.A1(net417),
    .A2(_02240_),
    .B1(_02476_),
    .B2(net3654),
    .Y(_02757_));
 sky130_fd_sc_hd__o21ai_2 _20345_ (.A1(_02665_),
    .A2(_02756_),
    .B1(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__xnor3_1 _20346_ (.A(_02752_),
    .B(_02753_),
    .C(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__xor3_1 _20347_ (.A(_02733_),
    .B(_02748_),
    .C(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__maj3_1 _20348_ (.A(_02653_),
    .B(_02667_),
    .C(_02668_),
    .X(_02761_));
 sky130_fd_sc_hd__maj3_1 _20349_ (.A(_02647_),
    .B(_02651_),
    .C(_02652_),
    .X(_02762_));
 sky130_fd_sc_hd__maj3_1 _20350_ (.A(_02673_),
    .B(_02674_),
    .C(_02675_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_8 _20351_ (.A0(_09243_),
    .A1(_10294_),
    .S(net3760),
    .X(_02764_));
 sky130_fd_sc_hd__nor2_2 _20352_ (.A(net3657),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_2 _20353_ (.A(net3661),
    .B(_02505_),
    .Y(_02766_));
 sky130_fd_sc_hd__nor2_2 _20354_ (.A(net3648),
    .B(_02680_),
    .Y(_02767_));
 sky130_fd_sc_hd__xnor3_1 _20355_ (.A(_02765_),
    .B(_02766_),
    .C(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__nor2_1 _20356_ (.A(net3653),
    .B(_02318_),
    .Y(_02769_));
 sky130_fd_sc_hd__nor2_1 _20357_ (.A(net446),
    .B(net3638),
    .Y(_02770_));
 sky130_fd_sc_hd__nor2_1 _20358_ (.A(_01693_),
    .B(net3635),
    .Y(_02771_));
 sky130_fd_sc_hd__xnor3_1 _20359_ (.A(_02769_),
    .B(_02770_),
    .C(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__xor3_1 _20360_ (.A(_02763_),
    .B(_02768_),
    .C(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__maj3_1 _20361_ (.A(_02672_),
    .B(_02676_),
    .C(_02682_),
    .X(_02774_));
 sky130_fd_sc_hd__xnor3_1 _20362_ (.A(_02762_),
    .B(_02773_),
    .C(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__xnor2_1 _20363_ (.A(_02761_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_2 _20364_ (.A(_02760_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__xnor3_1 _20365_ (.A(_02653_),
    .B(_02667_),
    .C(_02668_),
    .X(_02778_));
 sky130_fd_sc_hd__maj3_4 _20366_ (.A(_02778_),
    .B(_02685_),
    .C(_02687_),
    .X(_02779_));
 sky130_fd_sc_hd__nor2_4 _20367_ (.A(net3648),
    .B(_02764_),
    .Y(_02780_));
 sky130_fd_sc_hd__nor4_1 _20368_ (.A(net3657),
    .B(_01762_),
    .C(_02505_),
    .D(_02680_),
    .Y(_02781_));
 sky130_fd_sc_hd__o22ai_1 _20369_ (.A1(net3657),
    .A2(_02505_),
    .B1(_02680_),
    .B2(_01762_),
    .Y(_02782_));
 sky130_fd_sc_hd__o21ai_4 _20370_ (.A1(_02780_),
    .A2(_02781_),
    .B1(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__mux2i_4 _20371_ (.A0(net3696),
    .A1(_10474_),
    .S(net3759),
    .Y(_02784_));
 sky130_fd_sc_hd__or2_4 _20372_ (.A(_01762_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__xor2_1 _20373_ (.A(_02783_),
    .B(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__a21o_1 _20374_ (.A1(_02489_),
    .A2(_02565_),
    .B1(_02566_),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_1 _20375_ (.A(_02568_),
    .B(_02571_),
    .Y(_02788_));
 sky130_fd_sc_hd__maj3_1 _20376_ (.A(_02787_),
    .B(_02788_),
    .C(_02575_),
    .X(_02789_));
 sky130_fd_sc_hd__xor3_1 _20377_ (.A(_02672_),
    .B(_02676_),
    .C(_02682_),
    .X(_02790_));
 sky130_fd_sc_hd__maj3_1 _20378_ (.A(_02789_),
    .B(_02790_),
    .C(_02684_),
    .X(_02791_));
 sky130_fd_sc_hd__xnor2_1 _20379_ (.A(_02786_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__xor2_1 _20380_ (.A(_02779_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__xnor2_1 _20381_ (.A(_02777_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__xnor2_1 _20382_ (.A(_02669_),
    .B(_02687_),
    .Y(_02795_));
 sky130_fd_sc_hd__xnor2_1 _20383_ (.A(_02685_),
    .B(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_2 _20384_ (.A(_02510_),
    .B(_02780_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand3_1 _20385_ (.A(_02689_),
    .B(_02797_),
    .C(_02692_),
    .Y(_02798_));
 sky130_fd_sc_hd__or2_0 _20386_ (.A(_02689_),
    .B(_02692_),
    .X(_02799_));
 sky130_fd_sc_hd__inv_1 _20387_ (.A(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__nand3_2 _20388_ (.A(_02691_),
    .B(_02796_),
    .C(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__o21ai_0 _20389_ (.A1(_02689_),
    .A2(_02692_),
    .B1(_02797_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_2 _20390_ (.A(_02689_),
    .B(_02692_),
    .Y(_02803_));
 sky130_fd_sc_hd__a22o_4 _20391_ (.A1(_02796_),
    .A2(_02798_),
    .B1(_02802_),
    .B2(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__maj3_1 _20392_ (.A(_02689_),
    .B(_02688_),
    .C(_02692_),
    .X(_02805_));
 sky130_fd_sc_hd__o22a_1 _20393_ (.A1(_02688_),
    .A2(_02799_),
    .B1(_02805_),
    .B2(_02797_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _20394_ (.A0(_02804_),
    .A1(_02806_),
    .S(_02644_),
    .X(_02807_));
 sky130_fd_sc_hd__o211ai_1 _20395_ (.A1(_02796_),
    .A2(_02798_),
    .B1(_02801_),
    .C1(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_1 _20396_ (.A(_02794_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_2 _20397_ (.A(_02600_),
    .B(_02696_),
    .Y(_02810_));
 sky130_fd_sc_hd__and2_0 _20398_ (.A(_02602_),
    .B(_02696_),
    .X(_02811_));
 sky130_fd_sc_hd__a31oi_2 _20399_ (.A1(_02525_),
    .A2(_02600_),
    .A3(_02696_),
    .B1(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__o21ai_4 _20400_ (.A1(_02550_),
    .A2(_02810_),
    .B1(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__xor2_4 _20401_ (.A(net3509),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__nor2_1 _20402_ (.A(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B(_02000_),
    .Y(_02815_));
 sky130_fd_sc_hd__a21oi_4 _20403_ (.A1(_02000_),
    .A2(_02814_),
    .B1(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__mux2_8 _20404_ (.A0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A1(_02816_),
    .S(_08009_),
    .X(_02817_));
 sky130_fd_sc_hd__nand2_1 _20405_ (.A(net3513),
    .B(_02006_),
    .Y(_02818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_486 ();
 sky130_fd_sc_hd__mux2i_4 _20407_ (.A0(_02217_),
    .A1(_02198_),
    .S(net3559),
    .Y(_02820_));
 sky130_fd_sc_hd__o21ai_4 _20408_ (.A1(_02171_),
    .A2(_02820_),
    .B1(_02612_),
    .Y(_02821_));
 sky130_fd_sc_hd__o21ai_4 _20409_ (.A1(_02056_),
    .A2(_02179_),
    .B1(_02078_),
    .Y(_02822_));
 sky130_fd_sc_hd__nor2_1 _20410_ (.A(_02016_),
    .B(_02175_),
    .Y(_02823_));
 sky130_fd_sc_hd__mux2i_1 _20411_ (.A0(_02396_),
    .A1(_02392_),
    .S(net3558),
    .Y(_02824_));
 sky130_fd_sc_hd__nor2_1 _20412_ (.A(_02056_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__or3_4 _20413_ (.A(net3557),
    .B(_02823_),
    .C(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__o21ai_4 _20414_ (.A1(net3560),
    .A2(_02822_),
    .B1(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_485 ();
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(_09337_),
    .B(net3589),
    .Y(_02829_));
 sky130_fd_sc_hd__xor2_1 _20417_ (.A(_02133_),
    .B(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__o21ai_0 _20418_ (.A1(_09337_),
    .A2(net3589),
    .B1(_02137_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21oi_1 _20419_ (.A1(_02127_),
    .A2(_02830_),
    .B1(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a221oi_1 _20420_ (.A1(net3603),
    .A2(_02821_),
    .B1(_02827_),
    .B2(net3602),
    .C1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand3_1 _20421_ (.A(net3746),
    .B(_02818_),
    .C(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__o21ai_2 _20422_ (.A1(net3746),
    .A2(_02817_),
    .B1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand3_4 _20423_ (.A(_11233_),
    .B(_01655_),
    .C(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2_8 _20424_ (.A(_02730_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_484 ();
 sky130_fd_sc_hd__nand2_1 _20426_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .B(_02153_),
    .Y(_02839_));
 sky130_fd_sc_hd__o21ai_0 _20427_ (.A1(_02153_),
    .A2(_02837_),
    .B1(_02839_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2b_1 _20428_ (.A_N(net56),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02840_));
 sky130_fd_sc_hd__o21ai_2 _20429_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net51),
    .B1(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__mux2_1 _20430_ (.A0(net33),
    .A1(net42),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_02842_));
 sky130_fd_sc_hd__nor2_1 _20431_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a211oi_2 _20432_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_02841_),
    .B1(_02843_),
    .C1(_10656_),
    .Y(_02844_));
 sky130_fd_sc_hd__inv_1 _20433_ (.A(\load_store_unit_i.rdata_q[15] ),
    .Y(_02845_));
 sky130_fd_sc_hd__o21ai_0 _20434_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .B1(_02840_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_8 _20435_ (.A(_10656_),
    .B(_10666_),
    .Y(_02847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_483 ();
 sky130_fd_sc_hd__a221oi_1 _20437_ (.A1(_02845_),
    .A2(_02420_),
    .B1(_02846_),
    .B2(net3822),
    .C1(_02847_),
    .Y(_02849_));
 sky130_fd_sc_hd__o32ai_2 _20438_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(\load_store_unit_i.rdata_offset_q[0] ),
    .A3(net33),
    .B1(_02844_),
    .B2(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand3_4 _20439_ (.A(net3472),
    .B(_01669_),
    .C(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_482 ();
 sky130_fd_sc_hd__maj3_4 _20441_ (.A(_02765_),
    .B(_02766_),
    .C(_02767_),
    .X(_02853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_481 ();
 sky130_fd_sc_hd__or2_4 _20443_ (.A(net3648),
    .B(_02784_),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_8 _20444_ (.A0(net390),
    .A1(_10390_),
    .S(net3760),
    .X(_02856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_480 ();
 sky130_fd_sc_hd__a21oi_1 _20446_ (.A1(_02783_),
    .A2(_02856_),
    .B1(_01762_),
    .Y(_02858_));
 sky130_fd_sc_hd__mux2i_4 _20447_ (.A0(net390),
    .A1(_10390_),
    .S(net3760),
    .Y(_02859_));
 sky130_fd_sc_hd__nor2_1 _20448_ (.A(_02784_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__mux2_1 _20449_ (.A0(_02860_),
    .A1(_02859_),
    .S(_02783_),
    .X(_02861_));
 sky130_fd_sc_hd__o21bai_1 _20450_ (.A1(net3648),
    .A2(_02783_),
    .B1_N(_02784_),
    .Y(_02862_));
 sky130_fd_sc_hd__a22oi_1 _20451_ (.A1(net3648),
    .A2(_02861_),
    .B1(_02862_),
    .B2(_02859_),
    .Y(_02863_));
 sky130_fd_sc_hd__o22ai_1 _20452_ (.A1(_02855_),
    .A2(_02858_),
    .B1(_02863_),
    .B2(_01762_),
    .Y(_02864_));
 sky130_fd_sc_hd__xnor2_1 _20453_ (.A(_02853_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__nor2_1 _20454_ (.A(_02676_),
    .B(_02682_),
    .Y(_02866_));
 sky130_fd_sc_hd__a21oi_1 _20455_ (.A1(_02676_),
    .A2(_02682_),
    .B1(_02672_),
    .Y(_02867_));
 sky130_fd_sc_hd__o21ai_0 _20456_ (.A1(_02866_),
    .A2(_02867_),
    .B1(_02773_),
    .Y(_02868_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(_02762_),
    .B(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__o31a_1 _20458_ (.A1(_02773_),
    .A2(_02866_),
    .A3(_02867_),
    .B1(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__xnor2_1 _20459_ (.A(_02865_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__maj3_4 _20460_ (.A(_02733_),
    .B(_02748_),
    .C(_02759_),
    .X(_02872_));
 sky130_fd_sc_hd__maj3_1 _20461_ (.A(_02736_),
    .B(_02740_),
    .C(_02747_),
    .X(_02873_));
 sky130_fd_sc_hd__maj3_2 _20462_ (.A(_02743_),
    .B(_02745_),
    .C(_02746_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2i_1 _20463_ (.A0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .S(_10740_),
    .Y(_02875_));
 sky130_fd_sc_hd__o22ai_2 _20464_ (.A1(_10422_),
    .A2(net3757),
    .B1(_02875_),
    .B2(_01738_),
    .Y(_02876_));
 sky130_fd_sc_hd__mux2_8 _20465_ (.A0(net3697),
    .A1(_10415_),
    .S(_01685_),
    .X(_02877_));
 sky130_fd_sc_hd__nor2_1 _20466_ (.A(_01711_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nor2_1 _20467_ (.A(_01700_),
    .B(_02744_),
    .Y(_02879_));
 sky130_fd_sc_hd__xor3_1 _20468_ (.A(_02876_),
    .B(_02878_),
    .C(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__nor2_1 _20469_ (.A(net3658),
    .B(_02583_),
    .Y(_02881_));
 sky130_fd_sc_hd__nor2_1 _20470_ (.A(net3654),
    .B(_02655_),
    .Y(_02882_));
 sky130_fd_sc_hd__nor2_1 _20471_ (.A(net417),
    .B(_02476_),
    .Y(_02883_));
 sky130_fd_sc_hd__xnor3_1 _20472_ (.A(_02881_),
    .B(_02882_),
    .C(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__xnor3_1 _20473_ (.A(_02874_),
    .B(_02880_),
    .C(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__maj3_1 _20474_ (.A(_02737_),
    .B(_02738_),
    .C(_02739_),
    .X(_02886_));
 sky130_fd_sc_hd__nor2_1 _20475_ (.A(net3643),
    .B(_02334_),
    .Y(_02887_));
 sky130_fd_sc_hd__nor2_1 _20476_ (.A(net3646),
    .B(net3639),
    .Y(_02888_));
 sky130_fd_sc_hd__nor2_1 _20477_ (.A(net3647),
    .B(_02240_),
    .Y(_02889_));
 sky130_fd_sc_hd__xor3_1 _20478_ (.A(_02887_),
    .B(_02888_),
    .C(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__maj3_1 _20479_ (.A(_02749_),
    .B(_02750_),
    .C(_02751_),
    .X(_02891_));
 sky130_fd_sc_hd__xnor3_1 _20480_ (.A(_02886_),
    .B(_02890_),
    .C(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__xnor3_1 _20481_ (.A(_02873_),
    .B(_02885_),
    .C(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__maj3_1 _20482_ (.A(_02763_),
    .B(_02768_),
    .C(_02772_),
    .X(_02894_));
 sky130_fd_sc_hd__maj3_1 _20483_ (.A(_02769_),
    .B(_02770_),
    .C(_02771_),
    .X(_02895_));
 sky130_fd_sc_hd__nor2_1 _20484_ (.A(net3653),
    .B(net3635),
    .Y(_02896_));
 sky130_fd_sc_hd__nor2_1 _20485_ (.A(_01745_),
    .B(net3638),
    .Y(_02897_));
 sky130_fd_sc_hd__nor2_1 _20486_ (.A(net3650),
    .B(_02318_),
    .Y(_02898_));
 sky130_fd_sc_hd__xor3_1 _20487_ (.A(_02896_),
    .B(_02897_),
    .C(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__mux2i_4 _20488_ (.A0(_09149_),
    .A1(_02679_),
    .S(net3760),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _20489_ (.A(_01886_),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__nor2_2 _20490_ (.A(_01693_),
    .B(_02505_),
    .Y(_02902_));
 sky130_fd_sc_hd__nor2_2 _20491_ (.A(net3661),
    .B(_02764_),
    .Y(_02903_));
 sky130_fd_sc_hd__xnor3_1 _20492_ (.A(_02901_),
    .B(_02902_),
    .C(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__xnor3_1 _20493_ (.A(_02895_),
    .B(_02899_),
    .C(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__maj3_4 _20494_ (.A(_02752_),
    .B(_02753_),
    .C(_02758_),
    .X(_02906_));
 sky130_fd_sc_hd__xnor3_1 _20495_ (.A(_02894_),
    .B(_02905_),
    .C(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__xnor2_1 _20496_ (.A(_02893_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_1 _20497_ (.A(_02872_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__maj3_1 _20498_ (.A(_02760_),
    .B(_02761_),
    .C(_02775_),
    .X(_02910_));
 sky130_fd_sc_hd__xnor2_1 _20499_ (.A(_02909_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__xnor2_1 _20500_ (.A(_02871_),
    .B(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__inv_1 _20501_ (.A(_02779_),
    .Y(_02913_));
 sky130_fd_sc_hd__and2_4 _20502_ (.A(_02786_),
    .B(_02791_),
    .X(_02914_));
 sky130_fd_sc_hd__inv_1 _20503_ (.A(_02684_),
    .Y(_02915_));
 sky130_fd_sc_hd__xnor3_1 _20504_ (.A(_02787_),
    .B(_02572_),
    .C(_02575_),
    .X(_02916_));
 sky130_fd_sc_hd__a21o_1 _20505_ (.A1(_02335_),
    .A2(_02466_),
    .B1(_02467_),
    .X(_02917_));
 sky130_fd_sc_hd__xor3_1 _20506_ (.A(_02469_),
    .B(_02470_),
    .C(_02471_),
    .X(_02918_));
 sky130_fd_sc_hd__maj3_1 _20507_ (.A(_02917_),
    .B(_02918_),
    .C(_02480_),
    .X(_02919_));
 sky130_fd_sc_hd__maj3_1 _20508_ (.A(_02916_),
    .B(_02590_),
    .C(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__nor2_1 _20509_ (.A(_02669_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nor3_1 _20510_ (.A(_02789_),
    .B(_02790_),
    .C(_02684_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _20511_ (.A(_02669_),
    .B(_02920_),
    .Y(_02923_));
 sky130_fd_sc_hd__a32oi_1 _20512_ (.A1(_02683_),
    .A2(_02915_),
    .A3(_02921_),
    .B1(_02922_),
    .B2(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__o211ai_1 _20513_ (.A1(_02683_),
    .A2(_02915_),
    .B1(_02921_),
    .C1(_02671_),
    .Y(_02925_));
 sky130_fd_sc_hd__a21oi_1 _20514_ (.A1(_02924_),
    .A2(_02925_),
    .B1(_02786_),
    .Y(_02926_));
 sky130_fd_sc_hd__nor2_1 _20515_ (.A(_02779_),
    .B(_02792_),
    .Y(_02927_));
 sky130_fd_sc_hd__nor3_1 _20516_ (.A(net3542),
    .B(_02914_),
    .C(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__a311oi_1 _20517_ (.A1(_02913_),
    .A2(_02777_),
    .A3(_02914_),
    .B1(_02926_),
    .C1(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__xnor2_1 _20518_ (.A(_02912_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__maj3_1 _20519_ (.A(_02691_),
    .B(_02796_),
    .C(_02803_),
    .X(_02931_));
 sky130_fd_sc_hd__o21bai_1 _20520_ (.A1(_02800_),
    .A2(_02931_),
    .B1_N(_02794_),
    .Y(_02932_));
 sky130_fd_sc_hd__and2_4 _20521_ (.A(_02801_),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__xnor2_1 _20522_ (.A(_02930_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__nor2_1 _20523_ (.A(_02697_),
    .B(_02809_),
    .Y(_02935_));
 sky130_fd_sc_hd__nand2_2 _20524_ (.A(_02644_),
    .B(_02695_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _20525_ (.A(_02602_),
    .B(_02696_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand2_1 _20526_ (.A(_02801_),
    .B(_02804_),
    .Y(_02938_));
 sky130_fd_sc_hd__xnor2_1 _20527_ (.A(_02794_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__a21oi_1 _20528_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__a31oi_1 _20529_ (.A1(_02603_),
    .A2(_02640_),
    .A3(_02935_),
    .B1(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__xnor2_4 _20530_ (.A(net3508),
    .B(net3489),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _20531_ (.A(_02000_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__o21ai_4 _20532_ (.A1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A2(_02000_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .Y(_02945_));
 sky130_fd_sc_hd__o21ai_4 _20534_ (.A1(net3937),
    .A2(_02944_),
    .B1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _20535_ (.A(net3507),
    .B(_02006_),
    .Y(_02947_));
 sky130_fd_sc_hd__o21ai_2 _20536_ (.A1(_11012_),
    .A2(_02058_),
    .B1(_02055_),
    .Y(_02948_));
 sky130_fd_sc_hd__mux2_1 _20537_ (.A0(_02446_),
    .A1(_02448_),
    .S(net3558),
    .X(_02949_));
 sky130_fd_sc_hd__nand2_1 _20538_ (.A(net3559),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__o211ai_1 _20539_ (.A1(net3559),
    .A2(_02053_),
    .B1(_02950_),
    .C1(net3560),
    .Y(_02951_));
 sky130_fd_sc_hd__o21ai_2 _20540_ (.A1(net3560),
    .A2(_02948_),
    .B1(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__mux2i_2 _20541_ (.A0(_02076_),
    .A1(_02098_),
    .S(_02016_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_2 _20542_ (.A1(net3557),
    .A2(_02953_),
    .B1(_02612_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(_09278_),
    .B(net3590),
    .Y(_02955_));
 sky130_fd_sc_hd__xor2_1 _20544_ (.A(_02133_),
    .B(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__o21ai_0 _20545_ (.A1(_09278_),
    .A2(net3590),
    .B1(_02137_),
    .Y(_02957_));
 sky130_fd_sc_hd__a21oi_1 _20546_ (.A1(_02127_),
    .A2(_02956_),
    .B1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__a221oi_2 _20547_ (.A1(net3602),
    .A2(_02952_),
    .B1(_02954_),
    .B2(net3603),
    .C1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand3_1 _20548_ (.A(net3744),
    .B(_02947_),
    .C(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__o21ai_2 _20549_ (.A1(net3744),
    .A2(_02946_),
    .B1(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__nand3_4 _20550_ (.A(_11253_),
    .B(_01655_),
    .C(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__nand2_8 _20551_ (.A(_02851_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__nand2_1 _20554_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .B(_02153_),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_0 _20555_ (.A1(_02153_),
    .A2(_02963_),
    .B1(_02966_),
    .Y(_00521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__nand2_1 _20558_ (.A(net3506),
    .B(_02006_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _20559_ (.A(_09491_),
    .B(net3588),
    .Y(_02970_));
 sky130_fd_sc_hd__xor2_1 _20560_ (.A(_02133_),
    .B(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__o21ai_0 _20561_ (.A1(_09491_),
    .A2(net3588),
    .B1(_02137_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_1 _20562_ (.A1(_02127_),
    .A2(_02971_),
    .B1(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__a221oi_1 _20563_ (.A1(net3603),
    .A2(_02952_),
    .B1(_02954_),
    .B2(net3602),
    .C1(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__nand3_1 _20564_ (.A(net3746),
    .B(_02969_),
    .C(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__a21oi_1 _20565_ (.A1(net3640),
    .A2(net3645),
    .B1(_01979_),
    .Y(_02976_));
 sky130_fd_sc_hd__nor2_4 _20566_ (.A(_01980_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__o21ai_0 _20567_ (.A1(_02602_),
    .A2(_02696_),
    .B1(_02525_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_2 _20568_ (.A(_02810_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_2 _20569_ (.A1(_02547_),
    .A2(_02549_),
    .B1(_02812_),
    .Y(_02980_));
 sky130_fd_sc_hd__nor2_1 _20570_ (.A(_02809_),
    .B(_02934_),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2b_1 _20571_ (.A(_02804_),
    .B_N(_02794_),
    .Y(_02982_));
 sky130_fd_sc_hd__a211oi_2 _20572_ (.A1(_02936_),
    .A2(_02933_),
    .B1(_02982_),
    .C1(_02930_),
    .Y(_02983_));
 sky130_fd_sc_hd__a31oi_4 _20573_ (.A1(_02979_),
    .A2(_02980_),
    .A3(_02981_),
    .B1(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__a22oi_2 _20575_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B1(_10746_),
    .B2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .Y(_02986_));
 sky130_fd_sc_hd__nand2_8 _20576_ (.A(_13078_),
    .B(_01685_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand2b_2 _20577_ (.A_N(net432),
    .B(net3757),
    .Y(_02988_));
 sky130_fd_sc_hd__nand3_2 _20578_ (.A(_09489_),
    .B(_13078_),
    .C(_01685_),
    .Y(_02989_));
 sky130_fd_sc_hd__or3_4 _20579_ (.A(net471),
    .B(net3744),
    .C(_10390_),
    .X(_02990_));
 sky130_fd_sc_hd__xnor2_1 _20580_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__o22ai_1 _20581_ (.A1(_02987_),
    .A2(_02988_),
    .B1(_02991_),
    .B2(net3757),
    .Y(_02992_));
 sky130_fd_sc_hd__xor2_1 _20582_ (.A(_02986_),
    .B(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__nor2_1 _20584_ (.A(_01700_),
    .B(_02877_),
    .Y(_02995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__nor2_1 _20586_ (.A(net3658),
    .B(_02655_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_2 _20587_ (.A(net3655),
    .B(_02744_),
    .Y(_02998_));
 sky130_fd_sc_hd__xnor2_1 _20588_ (.A(_02997_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__xnor2_1 _20589_ (.A(_02995_),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__maj3_1 _20590_ (.A(_02876_),
    .B(_02878_),
    .C(_02879_),
    .X(_03001_));
 sky130_fd_sc_hd__xor3_1 _20591_ (.A(_02993_),
    .B(_03000_),
    .C(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__a21bo_1 _20592_ (.A1(_02874_),
    .A2(_02880_),
    .B1_N(_02884_),
    .X(_03003_));
 sky130_fd_sc_hd__o21ai_2 _20593_ (.A1(_02874_),
    .A2(_02880_),
    .B1(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__nor2_1 _20594_ (.A(net417),
    .B(net3634),
    .Y(_03005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__nor2_1 _20596_ (.A(net3647),
    .B(_02334_),
    .Y(_03007_));
 sky130_fd_sc_hd__nor2_1 _20597_ (.A(net3643),
    .B(_02476_),
    .Y(_03008_));
 sky130_fd_sc_hd__xnor2_1 _20598_ (.A(_03007_),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__xnor2_1 _20599_ (.A(_03005_),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__maj3_1 _20600_ (.A(_02881_),
    .B(_02882_),
    .C(_02883_),
    .X(_03011_));
 sky130_fd_sc_hd__maj3_1 _20601_ (.A(_02887_),
    .B(_02888_),
    .C(_02889_),
    .X(_03012_));
 sky130_fd_sc_hd__xor2_1 _20602_ (.A(_03011_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__xnor2_1 _20603_ (.A(_03010_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__xnor2_1 _20604_ (.A(_03004_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__xnor2_2 _20605_ (.A(_03002_),
    .B(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__maj3_2 _20606_ (.A(_02896_),
    .B(_02897_),
    .C(_02898_),
    .X(_03017_));
 sky130_fd_sc_hd__or2_4 _20607_ (.A(net3646),
    .B(_02240_),
    .X(_03018_));
 sky130_fd_sc_hd__nor2_1 _20608_ (.A(net3639),
    .B(net3638),
    .Y(_03019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__nor2_1 _20610_ (.A(_01745_),
    .B(net3636),
    .Y(_03021_));
 sky130_fd_sc_hd__xnor3_1 _20611_ (.A(_03018_),
    .B(_03019_),
    .C(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__nor2_1 _20612_ (.A(net3653),
    .B(_02505_),
    .Y(_03023_));
 sky130_fd_sc_hd__nor2_1 _20613_ (.A(net3650),
    .B(net3635),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_1 _20614_ (.A(_01693_),
    .B(_02764_),
    .Y(_03025_));
 sky130_fd_sc_hd__xnor3_1 _20615_ (.A(_03023_),
    .B(_03024_),
    .C(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__xor2_1 _20616_ (.A(_03022_),
    .B(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__xnor2_1 _20617_ (.A(_03017_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__maj3_2 _20618_ (.A(_02886_),
    .B(_02890_),
    .C(_02891_),
    .X(_03029_));
 sky130_fd_sc_hd__maj3_1 _20619_ (.A(_02895_),
    .B(_02899_),
    .C(_02904_),
    .X(_03030_));
 sky130_fd_sc_hd__xnor2_1 _20620_ (.A(_03029_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__xnor2_1 _20621_ (.A(_03028_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__nand2b_1 _20622_ (.A_N(_02892_),
    .B(_02885_),
    .Y(_03033_));
 sky130_fd_sc_hd__nor2b_1 _20623_ (.A(_02885_),
    .B_N(_02892_),
    .Y(_03034_));
 sky130_fd_sc_hd__a21oi_2 _20624_ (.A1(_02873_),
    .A2(_03033_),
    .B1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_1 _20625_ (.A(_03032_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__xnor2_2 _20626_ (.A(_03016_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__inv_1 _20627_ (.A(_02893_),
    .Y(_03038_));
 sky130_fd_sc_hd__maj3_4 _20628_ (.A(_03038_),
    .B(_02872_),
    .C(_02907_),
    .X(_03039_));
 sky130_fd_sc_hd__maj3_4 _20629_ (.A(_02894_),
    .B(_02905_),
    .C(_02906_),
    .X(_03040_));
 sky130_fd_sc_hd__nand2_1 _20630_ (.A(_02765_),
    .B(_02766_),
    .Y(_03041_));
 sky130_fd_sc_hd__maj3_1 _20631_ (.A(_02900_),
    .B(_02765_),
    .C(_02766_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _20632_ (.A0(_03041_),
    .A1(_03042_),
    .S(_01778_),
    .X(_03043_));
 sky130_fd_sc_hd__xnor2_1 _20633_ (.A(_02856_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__or3_4 _20634_ (.A(_02783_),
    .B(_02785_),
    .C(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__nor2_1 _20636_ (.A(net3657),
    .B(_02784_),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_2 _20637_ (.A(net3648),
    .B(_02856_),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_1 _20638_ (.A(net3661),
    .B(_02680_),
    .Y(_03049_));
 sky130_fd_sc_hd__xor2_1 _20639_ (.A(_03048_),
    .B(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__xnor2_1 _20640_ (.A(_03047_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__a22o_1 _20641_ (.A1(_01886_),
    .A2(_02900_),
    .B1(_02902_),
    .B2(_02903_),
    .X(_03052_));
 sky130_fd_sc_hd__o21ai_2 _20642_ (.A1(_02902_),
    .A2(_02903_),
    .B1(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__xor2_2 _20643_ (.A(_03051_),
    .B(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__nor2_1 _20644_ (.A(net3648),
    .B(_02784_),
    .Y(_03055_));
 sky130_fd_sc_hd__maj3_1 _20645_ (.A(_02853_),
    .B(_03055_),
    .C(_02859_),
    .X(_03056_));
 sky130_fd_sc_hd__and2_0 _20646_ (.A(_02853_),
    .B(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__nor3_4 _20647_ (.A(net471),
    .B(net3747),
    .C(_10390_),
    .Y(_03058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__nand2_2 _20649_ (.A(net3760),
    .B(_03058_),
    .Y(_03060_));
 sky130_fd_sc_hd__a211oi_1 _20650_ (.A1(_02853_),
    .A2(_03055_),
    .B1(_03060_),
    .C1(net3644),
    .Y(_03061_));
 sky130_fd_sc_hd__a221o_1 _20651_ (.A1(net3644),
    .A2(_03056_),
    .B1(_03057_),
    .B2(_03060_),
    .C1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__xor2_2 _20652_ (.A(_03054_),
    .B(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__xnor2_1 _20653_ (.A(_03045_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__xnor2_1 _20654_ (.A(_03040_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__xnor2_1 _20655_ (.A(_03039_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__xnor2_1 _20656_ (.A(_03037_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nor2_1 _20657_ (.A(_02865_),
    .B(_02870_),
    .Y(_03068_));
 sky130_fd_sc_hd__inv_1 _20658_ (.A(_02910_),
    .Y(_03069_));
 sky130_fd_sc_hd__maj3_1 _20659_ (.A(_02871_),
    .B(_02909_),
    .C(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__xnor2_1 _20660_ (.A(_03068_),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__xnor2_2 _20661_ (.A(_03067_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__nand2_1 _20662_ (.A(_02779_),
    .B(_02792_),
    .Y(_03073_));
 sky130_fd_sc_hd__o21ai_2 _20663_ (.A1(_02777_),
    .A2(_02927_),
    .B1(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _20664_ (.A(_02914_),
    .B(_02912_),
    .Y(_03075_));
 sky130_fd_sc_hd__nor2_1 _20665_ (.A(_02914_),
    .B(_02912_),
    .Y(_03076_));
 sky130_fd_sc_hd__a21oi_2 _20666_ (.A1(_03074_),
    .A2(_03075_),
    .B1(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__xnor2_1 _20667_ (.A(_03072_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__xnor2_2 _20668_ (.A(_02984_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_1 _20669_ (.A(_02000_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__o21ai_4 _20670_ (.A1(_02000_),
    .A2(_02977_),
    .B1(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand2_1 _20671_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .Y(_03082_));
 sky130_fd_sc_hd__o211ai_1 _20672_ (.A1(net3937),
    .A2(_03081_),
    .B1(_03082_),
    .C1(net3755),
    .Y(_03083_));
 sky130_fd_sc_hd__a21oi_2 _20673_ (.A1(_02975_),
    .A2(_03083_),
    .B1(net3738),
    .Y(_03084_));
 sky130_fd_sc_hd__a21oi_4 _20674_ (.A1(net3738),
    .A2(_11268_),
    .B1(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__a21boi_4 _20675_ (.A1(\load_store_unit_i.data_sign_ext_q ),
    .A2(_02844_),
    .B1_N(_01669_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux4_2 _20676_ (.A0(net34),
    .A1(net27),
    .A2(\load_store_unit_i.rdata_q[16] ),
    .A3(net57),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_01670_),
    .B(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nand3_1 _20678_ (.A(net3472),
    .B(_03086_),
    .C(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__o21ai_2 _20679_ (.A1(net3472),
    .A2(_03085_),
    .B1(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__nand2_1 _20681_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .B(_02153_),
    .Y(_03092_));
 sky130_fd_sc_hd__o21ai_0 _20682_ (.A1(_02153_),
    .A2(net3447),
    .B1(_03092_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand3_4 _20683_ (.A(net3946),
    .B(net3827),
    .C(net3945),
    .Y(_03093_));
 sky130_fd_sc_hd__nand3_4 _20684_ (.A(net3829),
    .B(net3828),
    .C(_02150_),
    .Y(_03094_));
 sky130_fd_sc_hd__nor2_4 _20685_ (.A(_03093_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__o21ai_0 _20687_ (.A1(_01802_),
    .A2(_01979_),
    .B1(net3645),
    .Y(_03097_));
 sky130_fd_sc_hd__a21oi_1 _20688_ (.A1(_01778_),
    .A2(_01979_),
    .B1(_01711_),
    .Y(_03098_));
 sky130_fd_sc_hd__nand3_1 _20689_ (.A(_01700_),
    .B(net3640),
    .C(_01979_),
    .Y(_03099_));
 sky130_fd_sc_hd__o21ai_0 _20690_ (.A1(_01700_),
    .A2(_01979_),
    .B1(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(net3649),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__o21ai_0 _20692_ (.A1(_01700_),
    .A2(_03098_),
    .B1(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__a22oi_1 _20693_ (.A1(_01971_),
    .A2(_03097_),
    .B1(_03102_),
    .B2(net3645),
    .Y(_03103_));
 sky130_fd_sc_hd__xor2_2 _20694_ (.A(_01969_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__nor2_1 _20695_ (.A(_02792_),
    .B(_02801_),
    .Y(_03105_));
 sky130_fd_sc_hd__o21ai_0 _20696_ (.A1(_02913_),
    .A2(net3542),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2b_1 _20697_ (.A_N(_02792_),
    .B(_02804_),
    .Y(_03107_));
 sky130_fd_sc_hd__nand2_1 _20698_ (.A(_02801_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nand3_1 _20699_ (.A(_02913_),
    .B(net3542),
    .C(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__nand2_1 _20700_ (.A(_03106_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand2b_1 _20701_ (.A_N(_03072_),
    .B(_03075_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _20702_ (.A(_02933_),
    .B(_03074_),
    .Y(_03112_));
 sky130_fd_sc_hd__maj3_1 _20703_ (.A(_02914_),
    .B(_02912_),
    .C(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__a22oi_1 _20704_ (.A1(_03110_),
    .A2(_03111_),
    .B1(_03113_),
    .B2(_03072_),
    .Y(_03114_));
 sky130_fd_sc_hd__o31ai_1 _20705_ (.A1(_02934_),
    .A2(_02941_),
    .A3(_03078_),
    .B1(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__inv_1 _20706_ (.A(_03068_),
    .Y(_03116_));
 sky130_fd_sc_hd__maj3_4 _20707_ (.A(_03116_),
    .B(_03070_),
    .C(_03067_),
    .X(_03117_));
 sky130_fd_sc_hd__inv_1 _20708_ (.A(_02993_),
    .Y(_03118_));
 sky130_fd_sc_hd__maj3_2 _20709_ (.A(_03118_),
    .B(_03000_),
    .C(_03001_),
    .X(_03119_));
 sky130_fd_sc_hd__nand2_4 _20710_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .Y(_03120_));
 sky130_fd_sc_hd__a21boi_4 _20711_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(_10746_),
    .B1_N(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__nor2_4 _20712_ (.A(_13098_),
    .B(_01677_),
    .Y(_03122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__xnor2_1 _20714_ (.A(net3712),
    .B(net268),
    .Y(_03124_));
 sky130_fd_sc_hd__xnor2_1 _20715_ (.A(net409),
    .B(_09489_),
    .Y(_03125_));
 sky130_fd_sc_hd__mux2i_2 _20716_ (.A0(_03124_),
    .A1(_03125_),
    .S(_01681_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _20717_ (.A(_03122_),
    .B(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__xor2_1 _20718_ (.A(_03121_),
    .B(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__maj3_1 _20720_ (.A(_02986_),
    .B(_02989_),
    .C(_02990_),
    .X(_03130_));
 sky130_fd_sc_hd__o32a_1 _20721_ (.A1(_02986_),
    .A2(_02987_),
    .A3(_02988_),
    .B1(_03130_),
    .B2(net3757),
    .X(_03131_));
 sky130_fd_sc_hd__nor2_1 _20722_ (.A(net3658),
    .B(_02744_),
    .Y(_03132_));
 sky130_fd_sc_hd__nor2_1 _20723_ (.A(net3655),
    .B(_02877_),
    .Y(_03133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__nor2_1 _20725_ (.A(net3656),
    .B(net3633),
    .Y(_03135_));
 sky130_fd_sc_hd__xnor3_1 _20726_ (.A(_03132_),
    .B(_03133_),
    .C(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__xor2_1 _20727_ (.A(_03131_),
    .B(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__xnor2_1 _20728_ (.A(_03128_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__nor2_1 _20730_ (.A(net3643),
    .B(net3634),
    .Y(_03140_));
 sky130_fd_sc_hd__mux2i_4 _20731_ (.A0(net400),
    .A1(net3682),
    .S(_01685_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2_1 _20732_ (.A(_01783_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__nor2_1 _20734_ (.A(net3647),
    .B(_02476_),
    .Y(_03144_));
 sky130_fd_sc_hd__xnor2_1 _20735_ (.A(_03142_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__xnor2_1 _20736_ (.A(_03140_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__maj3_2 _20737_ (.A(_03005_),
    .B(_03007_),
    .C(_03008_),
    .X(_03147_));
 sky130_fd_sc_hd__maj3_2 _20738_ (.A(_02995_),
    .B(_02997_),
    .C(_02998_),
    .X(_03148_));
 sky130_fd_sc_hd__xor2_1 _20739_ (.A(_03147_),
    .B(_03148_),
    .X(_03149_));
 sky130_fd_sc_hd__xnor2_1 _20740_ (.A(_03146_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__xor2_1 _20741_ (.A(_03138_),
    .B(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__xnor2_1 _20742_ (.A(_03119_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__o21ai_0 _20744_ (.A1(net3639),
    .A2(net3638),
    .B1(_03018_),
    .Y(_03154_));
 sky130_fd_sc_hd__nor3_1 _20745_ (.A(net3639),
    .B(net3638),
    .C(_03018_),
    .Y(_03155_));
 sky130_fd_sc_hd__a21oi_2 _20746_ (.A1(_03021_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand2_1 _20747_ (.A(_02243_),
    .B(_02320_),
    .Y(_03157_));
 sky130_fd_sc_hd__nor2_1 _20748_ (.A(net3638),
    .B(_02240_),
    .Y(_03158_));
 sky130_fd_sc_hd__nor2_1 _20749_ (.A(net3639),
    .B(_02318_),
    .Y(_03159_));
 sky130_fd_sc_hd__xnor3_1 _20750_ (.A(_03157_),
    .B(_03158_),
    .C(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__nor2_1 _20751_ (.A(net3653),
    .B(_02764_),
    .Y(_03161_));
 sky130_fd_sc_hd__nor2_1 _20752_ (.A(net3650),
    .B(_02505_),
    .Y(_03162_));
 sky130_fd_sc_hd__nor2_1 _20753_ (.A(_01693_),
    .B(_02680_),
    .Y(_03163_));
 sky130_fd_sc_hd__xnor3_1 _20754_ (.A(_03161_),
    .B(_03162_),
    .C(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_1 _20755_ (.A(_03160_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__xnor2_1 _20756_ (.A(_03156_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__maj3_1 _20757_ (.A(_03010_),
    .B(_03011_),
    .C(_03012_),
    .X(_03167_));
 sky130_fd_sc_hd__inv_1 _20758_ (.A(_03026_),
    .Y(_03168_));
 sky130_fd_sc_hd__maj3_1 _20759_ (.A(_03017_),
    .B(_03022_),
    .C(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__xnor3_1 _20760_ (.A(_03166_),
    .B(_03167_),
    .C(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__maj3_1 _20761_ (.A(_03004_),
    .B(_03002_),
    .C(_03014_),
    .X(_03171_));
 sky130_fd_sc_hd__nand2_1 _20762_ (.A(_03170_),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__or2_0 _20763_ (.A(_03170_),
    .B(_03171_),
    .X(_03173_));
 sky130_fd_sc_hd__nand2_1 _20764_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__xor2_1 _20765_ (.A(_03152_),
    .B(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__nand2_1 _20766_ (.A(_03032_),
    .B(_03035_),
    .Y(_03176_));
 sky130_fd_sc_hd__nor2_1 _20767_ (.A(_03032_),
    .B(_03035_),
    .Y(_03177_));
 sky130_fd_sc_hd__a21oi_2 _20768_ (.A1(_03016_),
    .A2(_03176_),
    .B1(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand3_1 _20769_ (.A(net3644),
    .B(_02855_),
    .C(_02859_),
    .Y(_03179_));
 sky130_fd_sc_hd__o21ai_0 _20770_ (.A1(_02855_),
    .A2(_02859_),
    .B1(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__nor2_4 _20771_ (.A(net3757),
    .B(_02990_),
    .Y(_03181_));
 sky130_fd_sc_hd__maj3_1 _20772_ (.A(_03054_),
    .B(_03057_),
    .C(_03181_),
    .X(_03182_));
 sky130_fd_sc_hd__a32o_4 _20773_ (.A1(_02853_),
    .A2(_03054_),
    .A3(_03180_),
    .B1(_03182_),
    .B2(_01762_),
    .X(_03183_));
 sky130_fd_sc_hd__nand2b_1 _20774_ (.A_N(_02785_),
    .B(_03048_),
    .Y(_03184_));
 sky130_fd_sc_hd__maj3_1 _20775_ (.A(_03051_),
    .B(_03053_),
    .C(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__nor2_1 _20776_ (.A(net3657),
    .B(_02856_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor2_1 _20777_ (.A(net3661),
    .B(_02784_),
    .Y(_03187_));
 sky130_fd_sc_hd__or4_4 _20778_ (.A(net471),
    .B(_08498_),
    .C(_10390_),
    .D(net3757),
    .X(_03188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__nor2_1 _20780_ (.A(_01778_),
    .B(_03188_),
    .Y(_03190_));
 sky130_fd_sc_hd__xnor2_1 _20781_ (.A(_03187_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_1 _20782_ (.A(_03186_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__maj3_1 _20783_ (.A(_03047_),
    .B(_03048_),
    .C(_03049_),
    .X(_03193_));
 sky130_fd_sc_hd__maj3_1 _20784_ (.A(_03023_),
    .B(_03024_),
    .C(_03025_),
    .X(_03194_));
 sky130_fd_sc_hd__xor2_1 _20785_ (.A(_03193_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__xnor2_1 _20786_ (.A(_03192_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xor2_1 _20787_ (.A(_03185_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__maj3_1 _20788_ (.A(_03028_),
    .B(_03029_),
    .C(_03030_),
    .X(_03198_));
 sky130_fd_sc_hd__xnor2_1 _20789_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_1 _20790_ (.A(_03183_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__xnor2_1 _20791_ (.A(_03178_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__xnor2_1 _20792_ (.A(_03175_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__nor2_2 _20793_ (.A(_03039_),
    .B(_03063_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_2 _20794_ (.A(_03039_),
    .B(_03063_),
    .Y(_03204_));
 sky130_fd_sc_hd__o21ai_0 _20795_ (.A1(_03045_),
    .A2(_03203_),
    .B1(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _20796_ (.A(_03037_),
    .B(_03040_),
    .Y(_03206_));
 sky130_fd_sc_hd__o211ai_1 _20797_ (.A1(_03037_),
    .A2(_03040_),
    .B1(_03203_),
    .C1(_03045_),
    .Y(_03207_));
 sky130_fd_sc_hd__nor2_1 _20798_ (.A(_03037_),
    .B(_03040_),
    .Y(_03208_));
 sky130_fd_sc_hd__a211oi_1 _20799_ (.A1(_03037_),
    .A2(_03040_),
    .B1(_03204_),
    .C1(_03045_),
    .Y(_03209_));
 sky130_fd_sc_hd__a21oi_1 _20800_ (.A1(_03205_),
    .A2(_03208_),
    .B1(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__o211ai_1 _20801_ (.A1(_03205_),
    .A2(_03206_),
    .B1(_03207_),
    .C1(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__xnor2_1 _20802_ (.A(_03202_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nor2_4 _20803_ (.A(_03117_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand2_2 _20804_ (.A(_03117_),
    .B(_03212_),
    .Y(_03214_));
 sky130_fd_sc_hd__nor2b_2 _20805_ (.A(_03213_),
    .B_N(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__xor2_2 _20806_ (.A(net3477),
    .B(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_2 _20807_ (.A(_02000_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__o21ai_4 _20808_ (.A1(_02000_),
    .A2(_03104_),
    .B1(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__mux2_4 _20809_ (.A0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A1(_03218_),
    .S(_08009_),
    .X(_03219_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(net3512),
    .B(_02006_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_1 _20811_ (.A(_09426_),
    .B(net3613),
    .Y(_03221_));
 sky130_fd_sc_hd__xor2_1 _20812_ (.A(_02133_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__o21ai_0 _20813_ (.A1(_09426_),
    .A2(net3613),
    .B1(_02137_),
    .Y(_03223_));
 sky130_fd_sc_hd__a21oi_1 _20814_ (.A1(_02127_),
    .A2(_03222_),
    .B1(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a221oi_1 _20815_ (.A1(net3602),
    .A2(_02821_),
    .B1(_02827_),
    .B2(net3603),
    .C1(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand3_2 _20816_ (.A(net3746),
    .B(_03220_),
    .C(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__o21ai_1 _20817_ (.A1(net3748),
    .A2(_03219_),
    .B1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__mux4_2 _20819_ (.A0(net35),
    .A1(net38),
    .A2(\load_store_unit_i.rdata_q[17] ),
    .A3(net58),
    .S0(net3822),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03229_));
 sky130_fd_sc_hd__nand2_1 _20820_ (.A(_01670_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__and3_4 _20821_ (.A(net3472),
    .B(_03086_),
    .C(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__a31oi_2 _20822_ (.A1(_11292_),
    .A2(net3469),
    .A3(_03227_),
    .B1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand2_1 _20823_ (.A(_03095_),
    .B(net3446),
    .Y(_03233_));
 sky130_fd_sc_hd__nand2_1 _20824_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .B(_02153_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _20825_ (.A(_03233_),
    .B(_03234_),
    .Y(_00523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__nand2_1 _20827_ (.A(_02419_),
    .B(net53),
    .Y(_03236_));
 sky130_fd_sc_hd__nand2_8 _20828_ (.A(net3822),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_03237_));
 sky130_fd_sc_hd__nand2_2 _20829_ (.A(_10656_),
    .B(\load_store_unit_i.data_type_q[1] ),
    .Y(_03238_));
 sky130_fd_sc_hd__a22oi_1 _20830_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net47),
    .B1(_03238_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _20831_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(net30),
    .Y(_03240_));
 sky130_fd_sc_hd__nor2b_1 _20832_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B_N(net39),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _20833_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__o21ai_0 _20834_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03240_),
    .B1(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__a221o_1 _20835_ (.A1(\load_store_unit_i.rdata_q[12] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[4] ),
    .C1(_02847_),
    .X(_03244_));
 sky130_fd_sc_hd__o21ai_0 _20836_ (.A1(_01670_),
    .A2(_03243_),
    .B1(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o221ai_1 _20837_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03236_),
    .B1(_03237_),
    .B2(_03239_),
    .C1(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__nand2_2 _20838_ (.A(_11629_),
    .B(net3469),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _20839_ (.A(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B(_02225_),
    .Y(_03248_));
 sky130_fd_sc_hd__xor2_1 _20840_ (.A(_01986_),
    .B(_01990_),
    .X(_03249_));
 sky130_fd_sc_hd__nand2_2 _20841_ (.A(_02000_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nand2_2 _20842_ (.A(_03248_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__mux2i_2 _20843_ (.A0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A1(_03251_),
    .S(_08009_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand2_1 _20844_ (.A(net3536),
    .B(_02006_),
    .Y(_03253_));
 sky130_fd_sc_hd__o21ai_2 _20845_ (.A1(net3557),
    .A2(_02445_),
    .B1(_02612_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _20846_ (.A(_02056_),
    .B(_02609_),
    .Y(_03255_));
 sky130_fd_sc_hd__nor2_1 _20847_ (.A(net3594),
    .B(net3603),
    .Y(_03256_));
 sky130_fd_sc_hd__a21oi_1 _20848_ (.A1(_10203_),
    .A2(net3603),
    .B1(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__nand2_1 _20849_ (.A(_10173_),
    .B(net3603),
    .Y(_03258_));
 sky130_fd_sc_hd__o21ai_1 _20850_ (.A1(net3600),
    .A2(net3603),
    .B1(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__mux2i_1 _20851_ (.A0(_03257_),
    .A1(_03259_),
    .S(net3619),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_1 _20852_ (.A(_10098_),
    .B(net3603),
    .Y(_03261_));
 sky130_fd_sc_hd__o21ai_1 _20853_ (.A1(net3601),
    .A2(net3603),
    .B1(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__mux2i_1 _20854_ (.A0(_08810_),
    .A1(_09986_),
    .S(net3603),
    .Y(_03263_));
 sky130_fd_sc_hd__mux2i_1 _20855_ (.A0(_03262_),
    .A1(_03263_),
    .S(net3619),
    .Y(_03264_));
 sky130_fd_sc_hd__mux2i_1 _20856_ (.A0(_03260_),
    .A1(_03264_),
    .S(net3578),
    .Y(_03265_));
 sky130_fd_sc_hd__mux2_1 _20857_ (.A0(_02116_),
    .A1(_03265_),
    .S(net3558),
    .X(_03266_));
 sky130_fd_sc_hd__nand2_2 _20858_ (.A(_02016_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__nor2_1 _20859_ (.A(net3560),
    .B(_02436_),
    .Y(_03268_));
 sky130_fd_sc_hd__a31o_4 _20860_ (.A1(net3560),
    .A2(_03255_),
    .A3(_03267_),
    .B1(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__nor2_1 _20861_ (.A(net3594),
    .B(_10547_),
    .Y(_03270_));
 sky130_fd_sc_hd__xnor2_1 _20862_ (.A(net3726),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__o21a_4 _20863_ (.A1(_10937_),
    .A2(_02135_),
    .B1(_02124_),
    .X(_03272_));
 sky130_fd_sc_hd__nor2_4 _20864_ (.A(_02129_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__a221oi_2 _20865_ (.A1(net3594),
    .A2(_10547_),
    .B1(_02127_),
    .B2(_03271_),
    .C1(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a221oi_4 _20866_ (.A1(net3603),
    .A2(_03254_),
    .B1(_03269_),
    .B2(net3602),
    .C1(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__and3_4 _20867_ (.A(net3747),
    .B(_03253_),
    .C(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__a21oi_4 _20868_ (.A1(net3756),
    .A2(_03252_),
    .B1(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__o22ai_2 _20869_ (.A1(net3469),
    .A2(_03246_),
    .B1(_03247_),
    .B2(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__nand2_8 _20871_ (.A(_10519_),
    .B(_02151_),
    .Y(_03280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 ();
 sky130_fd_sc_hd__nand2_1 _20874_ (.A(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .B(_03280_),
    .Y(_03283_));
 sky130_fd_sc_hd__o21ai_0 _20875_ (.A1(net3459),
    .A2(_03280_),
    .B1(_03283_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _20876_ (.A(_02419_),
    .B(net36),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _20877_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(\load_store_unit_i.rdata_q[18] ),
    .Y(_03285_));
 sky130_fd_sc_hd__and2_0 _20878_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(net28),
    .X(_03286_));
 sky130_fd_sc_hd__a211oi_1 _20879_ (.A1(_02419_),
    .A2(net49),
    .B1(_03286_),
    .C1(_02423_),
    .Y(_03287_));
 sky130_fd_sc_hd__a311oi_1 _20880_ (.A1(_02423_),
    .A2(_03284_),
    .A3(_03285_),
    .B1(_03287_),
    .C1(_02847_),
    .Y(_03288_));
 sky130_fd_sc_hd__nand2_8 _20881_ (.A(net3472),
    .B(_03086_),
    .Y(_03289_));
 sky130_fd_sc_hd__nand2_1 _20882_ (.A(_09663_),
    .B(_09622_),
    .Y(_03290_));
 sky130_fd_sc_hd__xor2_1 _20883_ (.A(_02133_),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__o21ai_0 _20884_ (.A1(_09663_),
    .A2(_09622_),
    .B1(_02137_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _20885_ (.A1(_02127_),
    .A2(_03291_),
    .B1(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__a221oi_1 _20886_ (.A1(net3603),
    .A2(_02713_),
    .B1(_02715_),
    .B2(net3602),
    .C1(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__o211ai_1 _20887_ (.A1(net3497),
    .A2(_02702_),
    .B1(_03294_),
    .C1(net3745),
    .Y(_03295_));
 sky130_fd_sc_hd__nor2_2 _20888_ (.A(_03072_),
    .B(_03077_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_2 _20889_ (.A(_03072_),
    .B(_03077_),
    .Y(_03297_));
 sky130_fd_sc_hd__o21ai_1 _20890_ (.A1(_02984_),
    .A2(_03296_),
    .B1(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__a21oi_2 _20891_ (.A1(_03214_),
    .A2(_03298_),
    .B1(_03213_),
    .Y(_03299_));
 sky130_fd_sc_hd__nor2_1 _20892_ (.A(_03131_),
    .B(_03136_),
    .Y(_03300_));
 sky130_fd_sc_hd__nand2_1 _20893_ (.A(_03131_),
    .B(_03136_),
    .Y(_03301_));
 sky130_fd_sc_hd__o21ai_2 _20894_ (.A1(_03128_),
    .A2(_03300_),
    .B1(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__nor2_2 _20895_ (.A(net3655),
    .B(_02987_),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _20896_ (.A(net3656),
    .B(_02744_),
    .Y(_03304_));
 sky130_fd_sc_hd__nor2_1 _20897_ (.A(net3658),
    .B(_02877_),
    .Y(_03305_));
 sky130_fd_sc_hd__xor3_1 _20898_ (.A(_03303_),
    .B(_03304_),
    .C(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__a2111oi_4 _20899_ (.A1(net432),
    .A2(net3757),
    .B1(_01677_),
    .C1(net387),
    .D1(_13098_),
    .Y(_03307_));
 sky130_fd_sc_hd__nor4_2 _20900_ (.A(_13098_),
    .B(_01698_),
    .C(net443),
    .D(_01677_),
    .Y(_03308_));
 sky130_fd_sc_hd__maj3_1 _20901_ (.A(_03121_),
    .B(_03307_),
    .C(net3627),
    .X(_03309_));
 sky130_fd_sc_hd__nor3_4 _20902_ (.A(_08498_),
    .B(_13076_),
    .C(_03120_),
    .Y(_03310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 ();
 sky130_fd_sc_hd__a21o_1 _20904_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_10746_),
    .B1(_03310_),
    .X(_03312_));
 sky130_fd_sc_hd__xnor2_1 _20905_ (.A(_03309_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__xnor2_1 _20906_ (.A(_03306_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 ();
 sky130_fd_sc_hd__o22ai_1 _20908_ (.A1(net3646),
    .A2(_02334_),
    .B1(_02476_),
    .B2(net3647),
    .Y(_03316_));
 sky130_fd_sc_hd__nor4_1 _20909_ (.A(net3647),
    .B(net3646),
    .C(_02334_),
    .D(_02476_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _20910_ (.A1(_03140_),
    .A2(_03316_),
    .B1(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__nor2_1 _20911_ (.A(net3647),
    .B(net3634),
    .Y(_03319_));
 sky130_fd_sc_hd__nor2_2 _20912_ (.A(net3641),
    .B(net3633),
    .Y(_03320_));
 sky130_fd_sc_hd__nor2_1 _20913_ (.A(net3646),
    .B(_02476_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor3_1 _20914_ (.A(_03319_),
    .B(_03320_),
    .C(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 ();
 sky130_fd_sc_hd__nor4_1 _20916_ (.A(net3658),
    .B(net3655),
    .C(_02744_),
    .D(_02877_),
    .Y(_03324_));
 sky130_fd_sc_hd__o22ai_1 _20917_ (.A1(net3658),
    .A2(_02744_),
    .B1(_02877_),
    .B2(net3655),
    .Y(_03325_));
 sky130_fd_sc_hd__o21ai_2 _20918_ (.A1(_03135_),
    .A2(_03324_),
    .B1(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__xnor3_1 _20919_ (.A(_03318_),
    .B(_03322_),
    .C(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__nand2_1 _20920_ (.A(_03314_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__or2_0 _20921_ (.A(_03314_),
    .B(_03327_),
    .X(_03329_));
 sky130_fd_sc_hd__nand2_1 _20922_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__xor2_1 _20923_ (.A(_03302_),
    .B(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 ();
 sky130_fd_sc_hd__o22ai_1 _20925_ (.A1(net3639),
    .A2(net3636),
    .B1(_02240_),
    .B2(net3638),
    .Y(_03333_));
 sky130_fd_sc_hd__nor4_1 _20926_ (.A(net3639),
    .B(net3638),
    .C(net3636),
    .D(_02240_),
    .Y(_03334_));
 sky130_fd_sc_hd__a31oi_1 _20927_ (.A1(_02243_),
    .A2(_02320_),
    .A3(_03333_),
    .B1(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__nor2_1 _20928_ (.A(net3639),
    .B(net3635),
    .Y(_03336_));
 sky130_fd_sc_hd__nor2_1 _20929_ (.A(net3638),
    .B(_02334_),
    .Y(_03337_));
 sky130_fd_sc_hd__nor2_1 _20930_ (.A(net3636),
    .B(_02240_),
    .Y(_03338_));
 sky130_fd_sc_hd__xnor3_1 _20931_ (.A(_03336_),
    .B(_03337_),
    .C(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__nor2_1 _20932_ (.A(net3653),
    .B(_02680_),
    .Y(_03340_));
 sky130_fd_sc_hd__nor2_1 _20933_ (.A(_01745_),
    .B(_02505_),
    .Y(_03341_));
 sky130_fd_sc_hd__nor2_1 _20934_ (.A(net3650),
    .B(_02764_),
    .Y(_03342_));
 sky130_fd_sc_hd__xnor3_1 _20935_ (.A(_03340_),
    .B(_03341_),
    .C(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__xor2_1 _20936_ (.A(_03339_),
    .B(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__xnor2_1 _20937_ (.A(_03335_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__inv_1 _20938_ (.A(_03164_),
    .Y(_03346_));
 sky130_fd_sc_hd__nor2_1 _20939_ (.A(_03160_),
    .B(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _20940_ (.A(_03160_),
    .B(_03346_),
    .Y(_03348_));
 sky130_fd_sc_hd__o21ai_2 _20941_ (.A1(_03156_),
    .A2(_03347_),
    .B1(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _20942_ (.A(_03147_),
    .B(_03148_),
    .Y(_03350_));
 sky130_fd_sc_hd__nor2_1 _20943_ (.A(_03147_),
    .B(_03148_),
    .Y(_03351_));
 sky130_fd_sc_hd__a21oi_1 _20944_ (.A1(_03146_),
    .A2(_03350_),
    .B1(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__xnor2_1 _20945_ (.A(_03349_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_1 _20946_ (.A(_03345_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nor2_1 _20947_ (.A(_03119_),
    .B(_03150_),
    .Y(_03355_));
 sky130_fd_sc_hd__nand2_1 _20948_ (.A(_03119_),
    .B(_03150_),
    .Y(_03356_));
 sky130_fd_sc_hd__o21ai_1 _20949_ (.A1(_03138_),
    .A2(_03355_),
    .B1(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__xor2_1 _20950_ (.A(_03354_),
    .B(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__xnor2_1 _20951_ (.A(_03331_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_2 _20952_ (.A(_03185_),
    .B(_03196_),
    .Y(_03360_));
 sky130_fd_sc_hd__maj3_1 _20953_ (.A(_03166_),
    .B(_03167_),
    .C(_03169_),
    .X(_03361_));
 sky130_fd_sc_hd__nand2b_2 _20954_ (.A_N(_02784_),
    .B(_01818_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_1 _20955_ (.A(_01815_),
    .B(_02859_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3_1 _20956_ (.A(net3760),
    .B(net3657),
    .C(_03058_),
    .Y(_03364_));
 sky130_fd_sc_hd__xor2_1 _20957_ (.A(_03363_),
    .B(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__xnor2_1 _20958_ (.A(_03362_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__maj3_1 _20959_ (.A(_03187_),
    .B(_03186_),
    .C(_03190_),
    .X(_03367_));
 sky130_fd_sc_hd__maj3_1 _20960_ (.A(_03161_),
    .B(_03162_),
    .C(_03163_),
    .X(_03368_));
 sky130_fd_sc_hd__xnor2_1 _20961_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__xnor2_1 _20962_ (.A(_03366_),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__maj3_1 _20963_ (.A(_03192_),
    .B(_03193_),
    .C(_03194_),
    .X(_03371_));
 sky130_fd_sc_hd__xor2_1 _20964_ (.A(_03370_),
    .B(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__xnor2_1 _20965_ (.A(_03361_),
    .B(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__xor2_1 _20966_ (.A(_03360_),
    .B(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__a21boi_0 _20967_ (.A1(_03152_),
    .A2(_03172_),
    .B1_N(_03173_),
    .Y(_03375_));
 sky130_fd_sc_hd__or2_4 _20968_ (.A(_03374_),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__nand2_1 _20969_ (.A(_03374_),
    .B(_03375_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _20970_ (.A(_03376_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xor2_1 _20971_ (.A(_03359_),
    .B(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__nor2_1 _20972_ (.A(_03178_),
    .B(_03200_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _20973_ (.A(_03178_),
    .B(_03200_),
    .Y(_03381_));
 sky130_fd_sc_hd__o21ai_2 _20974_ (.A1(_03175_),
    .A2(_03380_),
    .B1(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__maj3_2 _20975_ (.A(_03197_),
    .B(_03183_),
    .C(_03198_),
    .X(_03383_));
 sky130_fd_sc_hd__xnor2_1 _20976_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_1 _20977_ (.A(_03379_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__or2_0 _20978_ (.A(_03045_),
    .B(_03040_),
    .X(_03386_));
 sky130_fd_sc_hd__o211ai_1 _20979_ (.A1(_03202_),
    .A2(_03203_),
    .B1(_03386_),
    .C1(_03037_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _20980_ (.A(_03045_),
    .B(_03040_),
    .Y(_03388_));
 sky130_fd_sc_hd__a21oi_1 _20981_ (.A1(_03037_),
    .A2(_03204_),
    .B1(_03203_),
    .Y(_03389_));
 sky130_fd_sc_hd__nor2_1 _20982_ (.A(_03388_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__a21boi_0 _20983_ (.A1(_03204_),
    .A2(_03386_),
    .B1_N(_03388_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _20984_ (.A(_03389_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__o21ai_0 _20985_ (.A1(_03202_),
    .A2(_03390_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__and2_4 _20986_ (.A(_03387_),
    .B(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__nand2_2 _20987_ (.A(_03385_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__or2_4 _20988_ (.A(_03385_),
    .B(_03394_),
    .X(_03396_));
 sky130_fd_sc_hd__nand2_1 _20989_ (.A(_03395_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__xnor2_2 _20990_ (.A(_03299_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__xor2_1 _20991_ (.A(_01972_),
    .B(_01981_),
    .X(_03399_));
 sky130_fd_sc_hd__xor2_1 _20992_ (.A(_01926_),
    .B(_01954_),
    .X(_03400_));
 sky130_fd_sc_hd__xnor2_2 _20993_ (.A(_03399_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__nor2_1 _20994_ (.A(_02000_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__a21oi_4 _20995_ (.A1(_02000_),
    .A2(_03398_),
    .B1(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__mux2i_1 _20996_ (.A0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A1(_03403_),
    .S(_08009_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_4 _20997_ (.A(net3755),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__a21oi_4 _20998_ (.A1(_03295_),
    .A2(_03405_),
    .B1(net3738),
    .Y(_03406_));
 sky130_fd_sc_hd__a21oi_4 _20999_ (.A1(net3738),
    .A2(_11315_),
    .B1(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__o22ai_2 _21000_ (.A1(_03288_),
    .A2(_03289_),
    .B1(_03407_),
    .B2(net3472),
    .Y(_03408_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_450 ();
 sky130_fd_sc_hd__nand2_1 _21002_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .B(_02153_),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ai_0 _21003_ (.A1(_02153_),
    .A2(net3425),
    .B1(_03410_),
    .Y(_00525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_449 ();
 sky130_fd_sc_hd__nand3_1 _21005_ (.A(_01954_),
    .B(_01975_),
    .C(_01980_),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_1 _21006_ (.A(_01926_),
    .B(_01972_),
    .Y(_03413_));
 sky130_fd_sc_hd__a21oi_1 _21007_ (.A1(_01926_),
    .A2(_01972_),
    .B1(_01954_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_0 _21008_ (.A1(_03413_),
    .A2(_03414_),
    .B1(_01981_),
    .Y(_03415_));
 sky130_fd_sc_hd__or3_1 _21009_ (.A(_01926_),
    .B(_01954_),
    .C(_01972_),
    .X(_03416_));
 sky130_fd_sc_hd__o211ai_1 _21010_ (.A1(_01973_),
    .A2(_03412_),
    .B1(_03415_),
    .C1(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__xnor2_2 _21011_ (.A(_01965_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__inv_1 _21012_ (.A(_03396_),
    .Y(_03419_));
 sky130_fd_sc_hd__a21oi_1 _21013_ (.A1(net3476),
    .A2(_03214_),
    .B1(_03213_),
    .Y(_03420_));
 sky130_fd_sc_hd__o21ai_1 _21014_ (.A1(_03419_),
    .A2(_03420_),
    .B1(_03395_),
    .Y(_03421_));
 sky130_fd_sc_hd__nand2_2 _21015_ (.A(_03370_),
    .B(_03371_),
    .Y(_03422_));
 sky130_fd_sc_hd__maj3_1 _21016_ (.A(_03345_),
    .B(_03349_),
    .C(_03352_),
    .X(_03423_));
 sky130_fd_sc_hd__nor2_1 _21017_ (.A(net3653),
    .B(_02784_),
    .Y(_03424_));
 sky130_fd_sc_hd__nor2_1 _21018_ (.A(_01693_),
    .B(_02856_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor2_1 _21019_ (.A(_01815_),
    .B(_03188_),
    .Y(_03426_));
 sky130_fd_sc_hd__xor2_1 _21020_ (.A(_03425_),
    .B(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__xnor2_1 _21021_ (.A(_03424_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__maj3_2 _21022_ (.A(_03362_),
    .B(_03363_),
    .C(_03364_),
    .X(_03429_));
 sky130_fd_sc_hd__maj3_1 _21023_ (.A(_03340_),
    .B(_03341_),
    .C(_03342_),
    .X(_03430_));
 sky130_fd_sc_hd__xor2_1 _21024_ (.A(_03429_),
    .B(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__xnor2_1 _21025_ (.A(_03428_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__maj3_4 _21026_ (.A(_03366_),
    .B(_03367_),
    .C(_03368_),
    .X(_03433_));
 sky130_fd_sc_hd__xnor2_1 _21027_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _21028_ (.A(_03423_),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__or2_0 _21029_ (.A(_03423_),
    .B(_03434_),
    .X(_03436_));
 sky130_fd_sc_hd__nand2_1 _21030_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__xor2_1 _21031_ (.A(_03422_),
    .B(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__maj3_1 _21032_ (.A(_03331_),
    .B(_03354_),
    .C(_03357_),
    .X(_03439_));
 sky130_fd_sc_hd__nor2_2 _21033_ (.A(net3646),
    .B(net3634),
    .Y(_03440_));
 sky130_fd_sc_hd__nor2_1 _21034_ (.A(net3641),
    .B(_02744_),
    .Y(_03441_));
 sky130_fd_sc_hd__nor2_1 _21035_ (.A(net3647),
    .B(net3633),
    .Y(_03442_));
 sky130_fd_sc_hd__xor2_1 _21036_ (.A(_03441_),
    .B(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__xnor2_1 _21037_ (.A(_03440_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__maj3_4 _21038_ (.A(_03319_),
    .B(_03320_),
    .C(_03321_),
    .X(_03445_));
 sky130_fd_sc_hd__maj3_1 _21039_ (.A(_03303_),
    .B(_03304_),
    .C(_03305_),
    .X(_03446_));
 sky130_fd_sc_hd__xnor2_1 _21040_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__xnor2_1 _21041_ (.A(_03444_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_448 ();
 sky130_fd_sc_hd__nor2_2 _21043_ (.A(_01888_),
    .B(net3656),
    .Y(_03450_));
 sky130_fd_sc_hd__nand2_1 _21044_ (.A(net3656),
    .B(_01887_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand3_1 _21045_ (.A(_01890_),
    .B(net3655),
    .C(_03122_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21oi_1 _21046_ (.A1(_03451_),
    .A2(_03452_),
    .B1(net3658),
    .Y(_03453_));
 sky130_fd_sc_hd__a21oi_2 _21047_ (.A1(_03303_),
    .A2(_03450_),
    .B1(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _21048_ (.A(net3656),
    .B(_02877_),
    .Y(_03455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__a21oi_1 _21050_ (.A1(net3658),
    .A2(net3655),
    .B1(_02987_),
    .Y(_03457_));
 sky130_fd_sc_hd__o22ai_4 _21051_ (.A1(_02877_),
    .A2(_03454_),
    .B1(_03455_),
    .B2(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_8 _21052_ (.A(net3640),
    .B(_03122_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand2_8 _21053_ (.A(_01802_),
    .B(_03122_),
    .Y(_03460_));
 sky130_fd_sc_hd__nor2_2 _21054_ (.A(_03459_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_2 _21055_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_10746_),
    .B1(_03310_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _21056_ (.A(_03459_),
    .B(_03460_),
    .Y(_03463_));
 sky130_fd_sc_hd__o21ai_0 _21057_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a21oi_2 _21058_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_10746_),
    .B1(_03310_),
    .Y(_03465_));
 sky130_fd_sc_hd__xnor2_1 _21059_ (.A(_03464_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__xnor2_1 _21060_ (.A(_03458_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 ();
 sky130_fd_sc_hd__nand2_8 _21063_ (.A(_03459_),
    .B(net3627),
    .Y(_03470_));
 sky130_fd_sc_hd__nor3_4 _21064_ (.A(net3747),
    .B(_13076_),
    .C(_03120_),
    .Y(_03471_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 ();
 sky130_fd_sc_hd__a21o_4 _21066_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_10746_),
    .B1(_03471_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2i_1 _21067_ (.A0(_03306_),
    .A1(_03470_),
    .S(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 ();
 sky130_fd_sc_hd__nand3_1 _21069_ (.A(_03121_),
    .B(_03460_),
    .C(_03473_),
    .Y(_03476_));
 sky130_fd_sc_hd__o31ai_1 _21070_ (.A1(_03460_),
    .A2(_03306_),
    .A3(_03473_),
    .B1(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 ();
 sky130_fd_sc_hd__a21oi_1 _21072_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_10746_),
    .B1(_03471_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand3_1 _21073_ (.A(_03459_),
    .B(_03460_),
    .C(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__o31ai_1 _21074_ (.A1(_03461_),
    .A2(_03306_),
    .A3(_03479_),
    .B1(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__a221oi_2 _21075_ (.A1(_03121_),
    .A2(_03474_),
    .B1(_03477_),
    .B2(net3629),
    .C1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor3_1 _21076_ (.A(_03448_),
    .B(_03467_),
    .C(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__maj3_1 _21077_ (.A(_03336_),
    .B(_03337_),
    .C(_03338_),
    .X(_03484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 ();
 sky130_fd_sc_hd__nor2_1 _21079_ (.A(_01745_),
    .B(_02764_),
    .Y(_03486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 ();
 sky130_fd_sc_hd__nor2_1 _21081_ (.A(net3650),
    .B(_02680_),
    .Y(_03488_));
 sky130_fd_sc_hd__nor2_1 _21082_ (.A(net3639),
    .B(_02505_),
    .Y(_03489_));
 sky130_fd_sc_hd__xnor2_1 _21083_ (.A(_03488_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__xnor2_1 _21084_ (.A(_03486_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_02240_),
    .B(net3635),
    .Y(_03492_));
 sky130_fd_sc_hd__nor2_1 _21086_ (.A(net3638),
    .B(_02476_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_1 _21087_ (.A(_02270_),
    .B(_03141_),
    .Y(_03494_));
 sky130_fd_sc_hd__xor2_1 _21088_ (.A(_03493_),
    .B(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _21089_ (.A(_03492_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__xnor3_1 _21090_ (.A(_03484_),
    .B(_03491_),
    .C(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__maj3_1 _21091_ (.A(_03318_),
    .B(_03322_),
    .C(_03326_),
    .X(_03498_));
 sky130_fd_sc_hd__maj3_1 _21092_ (.A(_03335_),
    .B(_03339_),
    .C(_03343_),
    .X(_03499_));
 sky130_fd_sc_hd__nand2_1 _21093_ (.A(_03498_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__or2_0 _21094_ (.A(_03498_),
    .B(_03499_),
    .X(_03501_));
 sky130_fd_sc_hd__nand2_1 _21095_ (.A(_03500_),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__xnor2_1 _21096_ (.A(_03497_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__a21boi_1 _21097_ (.A1(_03302_),
    .A2(_03328_),
    .B1_N(_03329_),
    .Y(_03504_));
 sky130_fd_sc_hd__xnor2_1 _21098_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__xor2_1 _21099_ (.A(_03483_),
    .B(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__xnor2_1 _21100_ (.A(_03439_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _21101_ (.A(_03438_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__clkinv_1 _21102_ (.A(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__inv_1 _21103_ (.A(_03377_),
    .Y(_03510_));
 sky130_fd_sc_hd__o21ai_2 _21104_ (.A1(_03359_),
    .A2(_03510_),
    .B1(_03376_),
    .Y(_03511_));
 sky130_fd_sc_hd__maj3_1 _21105_ (.A(_03360_),
    .B(_03361_),
    .C(_03372_),
    .X(_03512_));
 sky130_fd_sc_hd__xnor2_1 _21106_ (.A(_03511_),
    .B(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__xnor2_1 _21107_ (.A(_03509_),
    .B(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__maj3_4 _21108_ (.A(_03382_),
    .B(_03379_),
    .C(_03383_),
    .X(_03515_));
 sky130_fd_sc_hd__xnor2_1 _21109_ (.A(net3488),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__xnor2_1 _21110_ (.A(net3468),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__nor2_2 _21111_ (.A(net3670),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__a21oi_4 _21112_ (.A1(net3670),
    .A2(_03418_),
    .B1(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__mux2i_4 _21113_ (.A0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A1(_03519_),
    .S(_08009_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _21114_ (.A(_09593_),
    .B(_09566_),
    .Y(_03521_));
 sky130_fd_sc_hd__xnor2_1 _21115_ (.A(_02133_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__o221ai_1 _21116_ (.A1(_09593_),
    .A2(_09566_),
    .B1(_02184_),
    .B2(_03522_),
    .C1(_02137_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _21117_ (.A(net3745),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__a21oi_1 _21118_ (.A1(net3602),
    .A2(_02617_),
    .B1(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__o21ai_0 _21119_ (.A1(_02020_),
    .A2(_02615_),
    .B1(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__a21oi_2 _21120_ (.A1(net160),
    .A2(_02006_),
    .B1(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__a21oi_4 _21121_ (.A1(net3755),
    .A2(_03520_),
    .B1(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__nand2_2 _21122_ (.A(net3738),
    .B(_11330_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21ai_4 _21123_ (.A1(net3738),
    .A2(_03528_),
    .B1(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__mux4_2 _21124_ (.A0(net37),
    .A1(net52),
    .A2(\load_store_unit_i.rdata_q[19] ),
    .A3(net29),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03531_));
 sky130_fd_sc_hd__a21oi_1 _21125_ (.A1(_01670_),
    .A2(_03531_),
    .B1(_03289_),
    .Y(_03532_));
 sky130_fd_sc_hd__a21oi_2 _21126_ (.A1(net3469),
    .A2(_03530_),
    .B1(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_439 ();
 sky130_fd_sc_hd__nand2_1 _21128_ (.A(_03095_),
    .B(net3416),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _21129_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .B(_02153_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _21130_ (.A(_03535_),
    .B(_03536_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _21131_ (.A(_03213_),
    .B(_03396_),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_2 _21132_ (.A(_03514_),
    .B(_03515_),
    .Y(_03538_));
 sky130_fd_sc_hd__a21oi_1 _21133_ (.A1(_03395_),
    .A2(_03537_),
    .B1(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _21134_ (.A(_03214_),
    .B(_03396_),
    .Y(_03540_));
 sky130_fd_sc_hd__a2111oi_0 _21135_ (.A1(_02984_),
    .A2(_03297_),
    .B1(_03296_),
    .C1(_03538_),
    .D1(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__a211o_4 _21136_ (.A1(net3488),
    .A2(_03515_),
    .B1(_03539_),
    .C1(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__maj3_4 _21137_ (.A(_03511_),
    .B(_03509_),
    .C(_03512_),
    .X(_03543_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_437 ();
 sky130_fd_sc_hd__a21o_4 _21140_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_10746_),
    .B1(_03310_),
    .X(_03546_));
 sky130_fd_sc_hd__nand3_1 _21141_ (.A(_03459_),
    .B(_03460_),
    .C(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_436 ();
 sky130_fd_sc_hd__nand2_1 _21143_ (.A(net3627),
    .B(_03465_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _21144_ (.A(net3629),
    .B(_03465_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_1 _21145_ (.A(net3627),
    .B(_03312_),
    .Y(_03551_));
 sky130_fd_sc_hd__a41o_1 _21146_ (.A1(_03547_),
    .A2(_03549_),
    .A3(_03550_),
    .A4(_03551_),
    .B1(_03458_),
    .X(_03552_));
 sky130_fd_sc_hd__nor4_1 _21147_ (.A(_03459_),
    .B(net3627),
    .C(_03462_),
    .D(_03546_),
    .Y(_03553_));
 sky130_fd_sc_hd__a21oi_1 _21148_ (.A1(_03461_),
    .A2(_03546_),
    .B1(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__o31a_1 _21149_ (.A1(_03462_),
    .A2(_03470_),
    .A3(_03546_),
    .B1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__o311ai_2 _21150_ (.A1(_03459_),
    .A2(_03462_),
    .A3(_03458_),
    .B1(_03552_),
    .C1(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__nor2_1 _21151_ (.A(net3641),
    .B(_02877_),
    .Y(_03557_));
 sky130_fd_sc_hd__nor2_1 _21152_ (.A(net3646),
    .B(net3633),
    .Y(_03558_));
 sky130_fd_sc_hd__nor2_1 _21153_ (.A(net3647),
    .B(_02744_),
    .Y(_03559_));
 sky130_fd_sc_hd__xor2_1 _21154_ (.A(_03558_),
    .B(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__xnor2_1 _21155_ (.A(_03557_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__maj3_1 _21156_ (.A(_03440_),
    .B(_03441_),
    .C(_03442_),
    .X(_03562_));
 sky130_fd_sc_hd__maj3_2 _21157_ (.A(net3658),
    .B(net3656),
    .C(net3655),
    .X(_03563_));
 sky130_fd_sc_hd__nand2b_4 _21158_ (.A_N(_03563_),
    .B(_03122_),
    .Y(_03564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_435 ();
 sky130_fd_sc_hd__xnor2_1 _21160_ (.A(_03562_),
    .B(_03564_),
    .Y(_03566_));
 sky130_fd_sc_hd__xnor2_1 _21161_ (.A(_03561_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__nor2_1 _21162_ (.A(net3658),
    .B(_01890_),
    .Y(_03568_));
 sky130_fd_sc_hd__o21ai_1 _21163_ (.A1(net3658),
    .A2(net3656),
    .B1(net3655),
    .Y(_03569_));
 sky130_fd_sc_hd__mux2i_4 _21164_ (.A0(net3697),
    .A1(_10415_),
    .S(_01685_),
    .Y(_03570_));
 sky130_fd_sc_hd__o311ai_4 _21165_ (.A1(net3655),
    .A2(_03450_),
    .A3(_03568_),
    .B1(_03569_),
    .C1(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand3_4 _21166_ (.A(net3658),
    .B(net3656),
    .C(net3655),
    .Y(_03572_));
 sky130_fd_sc_hd__a21bo_4 _21167_ (.A1(_03571_),
    .A2(_03572_),
    .B1_N(_03126_),
    .X(_03573_));
 sky130_fd_sc_hd__nand3b_1 _21168_ (.A_N(_03126_),
    .B(_03571_),
    .C(_03572_),
    .Y(_03574_));
 sky130_fd_sc_hd__a21oi_4 _21169_ (.A1(_03573_),
    .A2(_03574_),
    .B1(_02987_),
    .Y(_03575_));
 sky130_fd_sc_hd__a21oi_4 _21170_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(_10746_),
    .B1(_03471_),
    .Y(_03576_));
 sky130_fd_sc_hd__a21oi_1 _21171_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_10746_),
    .B1(_03471_),
    .Y(_03577_));
 sky130_fd_sc_hd__a21oi_1 _21172_ (.A1(net3627),
    .A2(_03546_),
    .B1(net3629),
    .Y(_03578_));
 sky130_fd_sc_hd__a21oi_1 _21173_ (.A1(_03460_),
    .A2(_03577_),
    .B1(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__xor2_1 _21174_ (.A(_03576_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__xnor2_1 _21175_ (.A(_03575_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__xor2_1 _21176_ (.A(_03567_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__xnor2_1 _21177_ (.A(_03556_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__nor2_1 _21178_ (.A(net3635),
    .B(_02334_),
    .Y(_03584_));
 sky130_fd_sc_hd__nor2_1 _21179_ (.A(net3638),
    .B(net3634),
    .Y(_03585_));
 sky130_fd_sc_hd__nor2_1 _21180_ (.A(net3636),
    .B(_02476_),
    .Y(_03586_));
 sky130_fd_sc_hd__xor2_1 _21181_ (.A(_03585_),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__xnor2_1 _21182_ (.A(_03584_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__inv_1 _21183_ (.A(_03494_),
    .Y(_03589_));
 sky130_fd_sc_hd__maj3_1 _21184_ (.A(_03492_),
    .B(_03493_),
    .C(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__nor2_1 _21185_ (.A(net3639),
    .B(_02764_),
    .Y(_03591_));
 sky130_fd_sc_hd__inv_1 _21186_ (.A(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _21187_ (.A(_02243_),
    .B(_02900_),
    .Y(_03593_));
 sky130_fd_sc_hd__or2_4 _21188_ (.A(_02240_),
    .B(_02505_),
    .X(_03594_));
 sky130_fd_sc_hd__xnor2_1 _21189_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__xnor2_1 _21190_ (.A(_03592_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__xnor2_1 _21191_ (.A(_03590_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__xnor2_1 _21192_ (.A(_03588_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__nand2_1 _21193_ (.A(_03445_),
    .B(_03446_),
    .Y(_03599_));
 sky130_fd_sc_hd__nor2_1 _21194_ (.A(_03445_),
    .B(_03446_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21oi_2 _21195_ (.A1(_03444_),
    .A2(_03599_),
    .B1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__maj3_1 _21196_ (.A(_03484_),
    .B(_03491_),
    .C(_03496_),
    .X(_03602_));
 sky130_fd_sc_hd__xnor2_1 _21197_ (.A(_03601_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_1 _21198_ (.A(_03598_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__inv_1 _21199_ (.A(_03482_),
    .Y(_03605_));
 sky130_fd_sc_hd__maj3_1 _21200_ (.A(_03448_),
    .B(_03467_),
    .C(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__xor2_1 _21201_ (.A(_03604_),
    .B(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__xnor2_1 _21202_ (.A(_03583_),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__inv_1 _21203_ (.A(_03504_),
    .Y(_03609_));
 sky130_fd_sc_hd__maj3_1 _21204_ (.A(_03483_),
    .B(_03503_),
    .C(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__inv_1 _21205_ (.A(_03500_),
    .Y(_03611_));
 sky130_fd_sc_hd__o21ai_1 _21206_ (.A1(_03497_),
    .A2(_03611_),
    .B1(_03501_),
    .Y(_03612_));
 sky130_fd_sc_hd__nor2b_2 _21207_ (.A(_03432_),
    .B_N(_03433_),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_1 _21208_ (.A(net3653),
    .B(_02856_),
    .Y(_03614_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(net3650),
    .B(_02784_),
    .Y(_03615_));
 sky130_fd_sc_hd__nor2_1 _21210_ (.A(_01818_),
    .B(_03188_),
    .Y(_03616_));
 sky130_fd_sc_hd__xnor2_1 _21211_ (.A(_03615_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__xnor2_1 _21212_ (.A(_03614_),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__maj3_1 _21213_ (.A(_03424_),
    .B(_03425_),
    .C(_03426_),
    .X(_03619_));
 sky130_fd_sc_hd__maj3_1 _21214_ (.A(_03486_),
    .B(_03488_),
    .C(_03489_),
    .X(_03620_));
 sky130_fd_sc_hd__xnor2_1 _21215_ (.A(_03619_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__xnor2_1 _21216_ (.A(_03618_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__inv_1 _21217_ (.A(_03430_),
    .Y(_03623_));
 sky130_fd_sc_hd__maj3_1 _21218_ (.A(_03429_),
    .B(_03428_),
    .C(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__xnor2_1 _21219_ (.A(_03622_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__xnor2_1 _21220_ (.A(_03613_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__xor2_1 _21221_ (.A(_03612_),
    .B(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_2 _21222_ (.A(_03610_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__or2_4 _21223_ (.A(_03610_),
    .B(_03627_),
    .X(_03629_));
 sky130_fd_sc_hd__nand2_1 _21224_ (.A(_03628_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__xor2_1 _21225_ (.A(_03608_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__inv_1 _21226_ (.A(_03506_),
    .Y(_03632_));
 sky130_fd_sc_hd__maj3_1 _21227_ (.A(_03439_),
    .B(_03632_),
    .C(_03438_),
    .X(_03633_));
 sky130_fd_sc_hd__a21boi_2 _21228_ (.A1(_03422_),
    .A2(_03435_),
    .B1_N(_03436_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_1 _21229_ (.A(_03633_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__xnor2_1 _21230_ (.A(_03631_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2_2 _21231_ (.A(_03543_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__or2_4 _21232_ (.A(_03543_),
    .B(_03636_),
    .X(_03638_));
 sky130_fd_sc_hd__nand2_1 _21233_ (.A(_03637_),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__xor2_1 _21234_ (.A(_03542_),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__nor2_2 _21235_ (.A(_02000_),
    .B(_03249_),
    .Y(_03641_));
 sky130_fd_sc_hd__a21oi_4 _21236_ (.A1(_02000_),
    .A2(_03640_),
    .B1(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__mux2i_2 _21237_ (.A0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A1(_03642_),
    .S(_08009_),
    .Y(_03643_));
 sky130_fd_sc_hd__nand2_1 _21238_ (.A(net3603),
    .B(_02453_),
    .Y(_03644_));
 sky130_fd_sc_hd__o21ai_2 _21239_ (.A1(_02057_),
    .A2(_02438_),
    .B1(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__inv_1 _21240_ (.A(_09797_),
    .Y(_03646_));
 sky130_fd_sc_hd__nand2_1 _21241_ (.A(_09790_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__xnor2_1 _21242_ (.A(_02133_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__o221ai_1 _21243_ (.A1(_09790_),
    .A2(_03646_),
    .B1(_02184_),
    .B2(_03648_),
    .C1(_02137_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_2 _21244_ (.A(net3746),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__a211oi_4 _21245_ (.A1(net161),
    .A2(_02006_),
    .B1(_03645_),
    .C1(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__a21oi_2 _21246_ (.A1(net3756),
    .A2(_03643_),
    .B1(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a211oi_1 _21247_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(\load_store_unit_i.rdata_q[20] ),
    .B1(_03241_),
    .C1(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_03653_));
 sky130_fd_sc_hd__a311o_1 _21248_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03240_),
    .A3(_03236_),
    .B1(_03653_),
    .C1(_02847_),
    .X(_03654_));
 sky130_fd_sc_hd__nand3_1 _21249_ (.A(net3472),
    .B(_03086_),
    .C(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o31ai_2 _21250_ (.A1(_11366_),
    .A2(net3472),
    .A3(_03652_),
    .B1(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_434 ();
 sky130_fd_sc_hd__nand2_1 _21252_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .B(_02153_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_0 _21253_ (.A1(_02153_),
    .A2(net3433),
    .B1(_03658_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _21254_ (.A(_09730_),
    .B(_09706_),
    .Y(_03659_));
 sky130_fd_sc_hd__xor2_1 _21255_ (.A(_03659_),
    .B(_02133_),
    .X(_03660_));
 sky130_fd_sc_hd__o21ai_0 _21256_ (.A1(_09730_),
    .A2(_09706_),
    .B1(_02137_),
    .Y(_03661_));
 sky130_fd_sc_hd__a21oi_1 _21257_ (.A1(_02127_),
    .A2(_03660_),
    .B1(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__a221oi_1 _21258_ (.A1(net3603),
    .A2(_02400_),
    .B1(_02405_),
    .B2(net3602),
    .C1(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__o211ai_1 _21259_ (.A1(net3496),
    .A2(_02702_),
    .B1(_03663_),
    .C1(net3745),
    .Y(_03664_));
 sky130_fd_sc_hd__nor2_1 _21260_ (.A(_08009_),
    .B(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .Y(_03665_));
 sky130_fd_sc_hd__a221oi_2 _21261_ (.A1(net3488),
    .A2(_03515_),
    .B1(_03543_),
    .B2(_03636_),
    .C1(_03421_),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _21262_ (.A(_03538_),
    .B(_03637_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand2_2 _21263_ (.A(_03638_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__nor2_1 _21264_ (.A(net3465),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__maj3_4 _21265_ (.A(_03633_),
    .B(_03631_),
    .C(_03634_),
    .X(_03670_));
 sky130_fd_sc_hd__maj3_1 _21266_ (.A(_03556_),
    .B(_03567_),
    .C(_03581_),
    .X(_03671_));
 sky130_fd_sc_hd__nor2_1 _21267_ (.A(net3641),
    .B(_02987_),
    .Y(_03672_));
 sky130_fd_sc_hd__nor2_1 _21268_ (.A(net3646),
    .B(_02744_),
    .Y(_03673_));
 sky130_fd_sc_hd__nor2_2 _21269_ (.A(net3647),
    .B(_02877_),
    .Y(_03674_));
 sky130_fd_sc_hd__xor2_1 _21270_ (.A(_03673_),
    .B(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__xnor2_1 _21271_ (.A(_03672_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__maj3_1 _21272_ (.A(_03557_),
    .B(_03558_),
    .C(_03559_),
    .X(_03677_));
 sky130_fd_sc_hd__xnor2_1 _21273_ (.A(_03564_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__xnor2_1 _21274_ (.A(_03676_),
    .B(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__nor2_1 _21275_ (.A(_03460_),
    .B(_03576_),
    .Y(_03680_));
 sky130_fd_sc_hd__nor2_4 _21276_ (.A(_01738_),
    .B(_10740_),
    .Y(_03681_));
 sky130_fd_sc_hd__a21oi_2 _21277_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(_03681_),
    .B1(_03471_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(_03460_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__o21ai_0 _21279_ (.A1(net3629),
    .A2(_03680_),
    .B1(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21oi_4 _21280_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_10746_),
    .B1(_03310_),
    .Y(_03685_));
 sky130_fd_sc_hd__xor2_1 _21281_ (.A(_03684_),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__xnor2_1 _21282_ (.A(_03575_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__xnor2_1 _21283_ (.A(_03679_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_432 ();
 sky130_fd_sc_hd__nand3_4 _21286_ (.A(_03122_),
    .B(_03571_),
    .C(_03572_),
    .Y(_03691_));
 sky130_fd_sc_hd__a21o_1 _21287_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_10746_),
    .B1(_03471_),
    .X(_03692_));
 sky130_fd_sc_hd__nor3_1 _21288_ (.A(net3627),
    .B(_03692_),
    .C(_03576_),
    .Y(_03693_));
 sky130_fd_sc_hd__a31oi_1 _21289_ (.A1(net3627),
    .A2(_03576_),
    .A3(_03691_),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_430 ();
 sky130_fd_sc_hd__nand2_4 _21292_ (.A(net3629),
    .B(net3627),
    .Y(_03697_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_429 ();
 sky130_fd_sc_hd__nand2_1 _21294_ (.A(_03692_),
    .B(_03576_),
    .Y(_03699_));
 sky130_fd_sc_hd__nand2_1 _21295_ (.A(net3627),
    .B(_03577_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand2_1 _21296_ (.A(_03460_),
    .B(_03576_),
    .Y(_03701_));
 sky130_fd_sc_hd__o21ai_0 _21297_ (.A1(_03576_),
    .A2(_03700_),
    .B1(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__a32oi_1 _21298_ (.A1(_03697_),
    .A2(_03691_),
    .A3(_03699_),
    .B1(_03702_),
    .B2(_03459_),
    .Y(_03703_));
 sky130_fd_sc_hd__o21ai_1 _21299_ (.A1(_03459_),
    .A2(_03694_),
    .B1(_03703_),
    .Y(_03704_));
 sky130_fd_sc_hd__xnor2_1 _21300_ (.A(_03688_),
    .B(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__inv_1 _21301_ (.A(_03561_),
    .Y(_03706_));
 sky130_fd_sc_hd__nor2_4 _21302_ (.A(_02987_),
    .B(_03563_),
    .Y(_03707_));
 sky130_fd_sc_hd__a21oi_1 _21303_ (.A1(_03706_),
    .A2(_03707_),
    .B1(_03562_),
    .Y(_03708_));
 sky130_fd_sc_hd__a21oi_2 _21304_ (.A1(_03561_),
    .A2(_03564_),
    .B1(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_1 _21305_ (.A(net3635),
    .B(_02476_),
    .Y(_03710_));
 sky130_fd_sc_hd__or2_4 _21306_ (.A(net3638),
    .B(net3633),
    .X(_03711_));
 sky130_fd_sc_hd__or2_4 _21307_ (.A(net3636),
    .B(net3634),
    .X(_03712_));
 sky130_fd_sc_hd__xnor2_1 _21308_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__xnor2_1 _21309_ (.A(_03710_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__maj3_1 _21310_ (.A(_03584_),
    .B(_03585_),
    .C(_03586_),
    .X(_03715_));
 sky130_fd_sc_hd__nor2_1 _21311_ (.A(net3639),
    .B(_02680_),
    .Y(_03716_));
 sky130_fd_sc_hd__nor2_1 _21312_ (.A(_02240_),
    .B(_02764_),
    .Y(_03717_));
 sky130_fd_sc_hd__nor2_1 _21313_ (.A(_02334_),
    .B(_02505_),
    .Y(_03718_));
 sky130_fd_sc_hd__xnor2_1 _21314_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__xnor2_1 _21315_ (.A(_03716_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__xor2_1 _21316_ (.A(_03715_),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__xnor2_1 _21317_ (.A(_03714_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _21318_ (.A(_03596_),
    .B(_03588_),
    .Y(_03723_));
 sky130_fd_sc_hd__nor2_1 _21319_ (.A(_03596_),
    .B(_03588_),
    .Y(_03724_));
 sky130_fd_sc_hd__a21o_1 _21320_ (.A1(_03590_),
    .A2(_03723_),
    .B1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__xor2_1 _21321_ (.A(_03722_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__xnor2_1 _21322_ (.A(_03709_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__xor2_1 _21323_ (.A(_03705_),
    .B(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__xnor2_1 _21324_ (.A(_03671_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__maj3_2 _21325_ (.A(_03601_),
    .B(_03598_),
    .C(_03602_),
    .X(_03730_));
 sky130_fd_sc_hd__inv_1 _21326_ (.A(_03624_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _21327_ (.A(_03622_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_1 _21328_ (.A(net3653),
    .B(_03181_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2b_1 _21329_ (.A_N(net3650),
    .B(_02859_),
    .Y(_03734_));
 sky130_fd_sc_hd__or2_4 _21330_ (.A(_01745_),
    .B(_02784_),
    .X(_03735_));
 sky130_fd_sc_hd__xnor2_1 _21331_ (.A(_03734_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__xnor2_1 _21332_ (.A(_03733_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__maj3_1 _21333_ (.A(_03614_),
    .B(_03615_),
    .C(_03616_),
    .X(_03738_));
 sky130_fd_sc_hd__maj3_2 _21334_ (.A(_03592_),
    .B(_03593_),
    .C(_03594_),
    .X(_03739_));
 sky130_fd_sc_hd__xnor2_1 _21335_ (.A(_03738_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__xnor2_1 _21336_ (.A(_03737_),
    .B(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__maj3_1 _21337_ (.A(_03619_),
    .B(_03618_),
    .C(_03620_),
    .X(_03742_));
 sky130_fd_sc_hd__xor2_1 _21338_ (.A(_03741_),
    .B(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__xnor2_1 _21339_ (.A(_03732_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__xnor2_1 _21340_ (.A(_03730_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__inv_1 _21341_ (.A(_03604_),
    .Y(_03746_));
 sky130_fd_sc_hd__maj3_1 _21342_ (.A(_03583_),
    .B(_03746_),
    .C(_03606_),
    .X(_03747_));
 sky130_fd_sc_hd__xnor2_1 _21343_ (.A(_03745_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__xnor2_1 _21344_ (.A(_03729_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2_2 _21345_ (.A(_03608_),
    .B(_03629_),
    .Y(_03750_));
 sky130_fd_sc_hd__maj3_1 _21346_ (.A(_03613_),
    .B(_03612_),
    .C(_03625_),
    .X(_03751_));
 sky130_fd_sc_hd__a21o_4 _21347_ (.A1(_03628_),
    .A2(_03750_),
    .B1(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__nand3_2 _21348_ (.A(_03628_),
    .B(_03751_),
    .C(_03750_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand2_1 _21349_ (.A(_03752_),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__xor2_1 _21350_ (.A(_03749_),
    .B(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__nor2_2 _21351_ (.A(_03670_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_2 _21352_ (.A(_03670_),
    .B(_03755_),
    .Y(_03757_));
 sky130_fd_sc_hd__inv_1 _21353_ (.A(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__nor2_1 _21354_ (.A(_03756_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__xor2_1 _21355_ (.A(_03669_),
    .B(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_1 _21356_ (.A(_01950_),
    .B(_01951_),
    .Y(_03761_));
 sky130_fd_sc_hd__xnor2_1 _21357_ (.A(_01952_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__nor2_1 _21358_ (.A(_01986_),
    .B(_01990_),
    .Y(_03763_));
 sky130_fd_sc_hd__xnor2_2 _21359_ (.A(_03762_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__nor2_1 _21360_ (.A(_02000_),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__a211oi_2 _21361_ (.A1(_02000_),
    .A2(_03760_),
    .B1(_03765_),
    .C1(net3937),
    .Y(_03766_));
 sky130_fd_sc_hd__o21ai_2 _21362_ (.A1(_03665_),
    .A2(_03766_),
    .B1(net3756),
    .Y(_03767_));
 sky130_fd_sc_hd__a21oi_4 _21363_ (.A1(_03664_),
    .A2(_03767_),
    .B1(net3738),
    .Y(_03768_));
 sky130_fd_sc_hd__a21oi_1 _21364_ (.A1(net3738),
    .A2(_11388_),
    .B1(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand2_2 _21365_ (.A(_02419_),
    .B(net54),
    .Y(_03770_));
 sky130_fd_sc_hd__nand2_1 _21366_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(net31),
    .Y(_03771_));
 sky130_fd_sc_hd__nor2b_1 _21367_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B_N(net40),
    .Y(_03772_));
 sky130_fd_sc_hd__a211oi_1 _21368_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(\load_store_unit_i.rdata_q[21] ),
    .B1(_03772_),
    .C1(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_03773_));
 sky130_fd_sc_hd__a311oi_1 _21369_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03770_),
    .A3(_03771_),
    .B1(_03773_),
    .C1(_02847_),
    .Y(_03774_));
 sky130_fd_sc_hd__o22ai_2 _21370_ (.A1(net3472),
    .A2(_03769_),
    .B1(_03774_),
    .B2(_03289_),
    .Y(_03775_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 ();
 sky130_fd_sc_hd__nand2_1 _21372_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .B(_02153_),
    .Y(_03777_));
 sky130_fd_sc_hd__o21ai_0 _21373_ (.A1(_02153_),
    .A2(net3413),
    .B1(_03777_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _21374_ (.A(_03637_),
    .B(_03757_),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_1 _21375_ (.A(_03542_),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nor2_1 _21376_ (.A(_03638_),
    .B(_03758_),
    .Y(_03780_));
 sky130_fd_sc_hd__nor3_1 _21377_ (.A(_03756_),
    .B(_03779_),
    .C(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_2 _21378_ (.A(_03749_),
    .B(_03753_),
    .Y(_03782_));
 sky130_fd_sc_hd__maj3_1 _21379_ (.A(_03671_),
    .B(_03705_),
    .C(_03727_),
    .X(_03783_));
 sky130_fd_sc_hd__xnor2_1 _21380_ (.A(net3641),
    .B(_01780_),
    .Y(_03784_));
 sky130_fd_sc_hd__a211oi_2 _21381_ (.A1(net3630),
    .A2(_03784_),
    .B1(net3646),
    .C1(_02877_),
    .Y(_03785_));
 sky130_fd_sc_hd__and3_4 _21382_ (.A(net3646),
    .B(net3630),
    .C(_03784_),
    .X(_03786_));
 sky130_fd_sc_hd__nor2_2 _21383_ (.A(_03785_),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__maj3_4 _21384_ (.A(_03672_),
    .B(_03673_),
    .C(_03674_),
    .X(_03788_));
 sky130_fd_sc_hd__xnor2_1 _21385_ (.A(_03707_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__xnor2_1 _21386_ (.A(_03787_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__inv_2 _21387_ (.A(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__a21o_4 _21388_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_03681_),
    .B1(_03471_),
    .X(_03792_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 ();
 sky130_fd_sc_hd__a21oi_1 _21390_ (.A1(net3627),
    .A2(_03792_),
    .B1(net3629),
    .Y(_03794_));
 sky130_fd_sc_hd__a21oi_1 _21391_ (.A1(_03460_),
    .A2(_03685_),
    .B1(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__a21o_4 _21392_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_03681_),
    .B1(_03471_),
    .X(_03796_));
 sky130_fd_sc_hd__xnor2_1 _21393_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__xnor2_1 _21394_ (.A(_03575_),
    .B(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__xnor2_1 _21395_ (.A(_03791_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__nand2_4 _21396_ (.A(_03697_),
    .B(_03691_),
    .Y(_03800_));
 sky130_fd_sc_hd__nor2_1 _21397_ (.A(_03682_),
    .B(_03792_),
    .Y(_03801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 ();
 sky130_fd_sc_hd__and3_4 _21399_ (.A(_03122_),
    .B(_03571_),
    .C(_03572_),
    .X(_03803_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 ();
 sky130_fd_sc_hd__nand3_1 _21401_ (.A(_03460_),
    .B(_03682_),
    .C(_03792_),
    .Y(_03805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_424 ();
 sky130_fd_sc_hd__o311ai_0 _21403_ (.A1(_03460_),
    .A2(_03792_),
    .A3(_03803_),
    .B1(_03805_),
    .C1(net3629),
    .Y(_03807_));
 sky130_fd_sc_hd__nand3_1 _21404_ (.A(net3627),
    .B(_03682_),
    .C(_03792_),
    .Y(_03808_));
 sky130_fd_sc_hd__o211ai_1 _21405_ (.A1(net3627),
    .A2(_03792_),
    .B1(_03808_),
    .C1(_03459_),
    .Y(_03809_));
 sky130_fd_sc_hd__a2bb2oi_2 _21406_ (.A1_N(_03800_),
    .A2_N(_03801_),
    .B1(_03807_),
    .B2(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__xor2_1 _21407_ (.A(_03799_),
    .B(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__inv_1 _21408_ (.A(_03676_),
    .Y(_03812_));
 sky130_fd_sc_hd__maj3_4 _21409_ (.A(_03707_),
    .B(_03812_),
    .C(_03677_),
    .X(_03813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_423 ();
 sky130_fd_sc_hd__nor2_1 _21411_ (.A(net3638),
    .B(_02744_),
    .Y(_03815_));
 sky130_fd_sc_hd__nor2_1 _21412_ (.A(net3635),
    .B(net3634),
    .Y(_03816_));
 sky130_fd_sc_hd__nor2_1 _21413_ (.A(net3636),
    .B(net3633),
    .Y(_03817_));
 sky130_fd_sc_hd__xor2_1 _21414_ (.A(_03816_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__xnor2_1 _21415_ (.A(_03815_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__inv_1 _21416_ (.A(_03710_),
    .Y(_03820_));
 sky130_fd_sc_hd__maj3_1 _21417_ (.A(_03820_),
    .B(_03711_),
    .C(_03712_),
    .X(_03821_));
 sky130_fd_sc_hd__nor2_1 _21418_ (.A(_02334_),
    .B(_02764_),
    .Y(_03822_));
 sky130_fd_sc_hd__nor2_1 _21419_ (.A(_02240_),
    .B(_02680_),
    .Y(_03823_));
 sky130_fd_sc_hd__nor2_1 _21420_ (.A(_02476_),
    .B(_02505_),
    .Y(_03824_));
 sky130_fd_sc_hd__xor2_1 _21421_ (.A(_03823_),
    .B(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__xnor2_1 _21422_ (.A(_03822_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__xor2_1 _21423_ (.A(_03821_),
    .B(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__xnor2_1 _21424_ (.A(_03819_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__maj3_1 _21425_ (.A(_03715_),
    .B(_03714_),
    .C(_03720_),
    .X(_03829_));
 sky130_fd_sc_hd__xor2_1 _21426_ (.A(_03828_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__xnor2_1 _21427_ (.A(_03813_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_422 ();
 sky130_fd_sc_hd__a21oi_2 _21429_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_10746_),
    .B1(_03471_),
    .Y(_03833_));
 sky130_fd_sc_hd__nor2_1 _21430_ (.A(net3627),
    .B(_03577_),
    .Y(_03834_));
 sky130_fd_sc_hd__a21oi_1 _21431_ (.A1(_03459_),
    .A2(_03700_),
    .B1(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__nor2_1 _21432_ (.A(net3627),
    .B(_03699_),
    .Y(_03836_));
 sky130_fd_sc_hd__o21ai_0 _21433_ (.A1(_03680_),
    .A2(_03836_),
    .B1(net3629),
    .Y(_03837_));
 sky130_fd_sc_hd__o21ai_0 _21434_ (.A1(_03470_),
    .A2(_03699_),
    .B1(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_1 _21435_ (.A(_03691_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__o31ai_1 _21436_ (.A1(_03576_),
    .A2(_03691_),
    .A3(_03835_),
    .B1(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__maj3_1 _21437_ (.A(_03576_),
    .B(_03803_),
    .C(_03835_),
    .X(_03841_));
 sky130_fd_sc_hd__xnor2_1 _21438_ (.A(_03833_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__and2_0 _21439_ (.A(_03679_),
    .B(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _21440_ (.A(net3627),
    .B(_03682_),
    .Y(_03844_));
 sky130_fd_sc_hd__o21ai_0 _21441_ (.A1(net3627),
    .A2(_03682_),
    .B1(net3629),
    .Y(_03845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_421 ();
 sky130_fd_sc_hd__a211oi_1 _21443_ (.A1(_03844_),
    .A2(_03845_),
    .B1(_03685_),
    .C1(_03691_),
    .Y(_03847_));
 sky130_fd_sc_hd__a211oi_2 _21444_ (.A1(_03833_),
    .A2(_03840_),
    .B1(_03843_),
    .C1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__xnor2_1 _21445_ (.A(_03831_),
    .B(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__xnor2_1 _21446_ (.A(_03811_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__inv_1 _21447_ (.A(_03722_),
    .Y(_03851_));
 sky130_fd_sc_hd__maj3_1 _21448_ (.A(_03851_),
    .B(_03709_),
    .C(_03725_),
    .X(_03852_));
 sky130_fd_sc_hd__nand2_1 _21449_ (.A(_03741_),
    .B(_03742_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _21450_ (.A(_03737_),
    .B(_03739_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand2_1 _21451_ (.A(_03738_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__o21ai_2 _21452_ (.A1(_03737_),
    .A2(_03739_),
    .B1(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_420 ();
 sky130_fd_sc_hd__or2_4 _21454_ (.A(net3639),
    .B(net3632),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_1 _21455_ (.A(_02243_),
    .B(_02859_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _21456_ (.A(net3650),
    .B(_03181_),
    .Y(_03860_));
 sky130_fd_sc_hd__xnor2_1 _21457_ (.A(_03859_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__xnor2_1 _21458_ (.A(_03858_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__maj3_1 _21459_ (.A(_03734_),
    .B(_03735_),
    .C(_03733_),
    .X(_03863_));
 sky130_fd_sc_hd__maj3_1 _21460_ (.A(_03717_),
    .B(_03716_),
    .C(_03718_),
    .X(_03864_));
 sky130_fd_sc_hd__inv_1 _21461_ (.A(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xnor2_1 _21462_ (.A(_03863_),
    .B(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__xnor2_1 _21463_ (.A(_03862_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__xnor2_1 _21464_ (.A(_03856_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_1 _21465_ (.A(_03853_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__xnor2_1 _21466_ (.A(_03852_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__xnor2_1 _21467_ (.A(_03850_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__xnor2_1 _21468_ (.A(_03783_),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _21469_ (.A(_03730_),
    .B(_03743_),
    .Y(_03873_));
 sky130_fd_sc_hd__nor2_1 _21470_ (.A(_03730_),
    .B(_03743_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21oi_1 _21471_ (.A1(_03732_),
    .A2(_03873_),
    .B1(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__inv_1 _21472_ (.A(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__maj3_1 _21473_ (.A(_03729_),
    .B(_03745_),
    .C(_03747_),
    .X(_03877_));
 sky130_fd_sc_hd__xnor2_1 _21474_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_1 _21475_ (.A(_03872_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__a21oi_2 _21476_ (.A1(_03752_),
    .A2(_03782_),
    .B1(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand3_2 _21477_ (.A(_03752_),
    .B(_03782_),
    .C(_03879_),
    .Y(_03881_));
 sky130_fd_sc_hd__nor2b_1 _21478_ (.A(_03880_),
    .B_N(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__xnor2_1 _21479_ (.A(_03781_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__or3_1 _21480_ (.A(net3544),
    .B(_01953_),
    .C(_01991_),
    .X(_03884_));
 sky130_fd_sc_hd__and2_4 _21481_ (.A(net3531),
    .B(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(_02000_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__a21oi_4 _21483_ (.A1(_02000_),
    .A2(_03883_),
    .B1(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__mux2i_2 _21484_ (.A0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A1(_03887_),
    .S(_08009_),
    .Y(_03888_));
 sky130_fd_sc_hd__nor2_1 _21485_ (.A(net436),
    .B(_09866_),
    .Y(_03889_));
 sky130_fd_sc_hd__xor2_1 _21486_ (.A(_02133_),
    .B(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__nand2_1 _21487_ (.A(net436),
    .B(_09866_),
    .Y(_03891_));
 sky130_fd_sc_hd__o211ai_1 _21488_ (.A1(_02184_),
    .A2(_03890_),
    .B1(_03891_),
    .C1(_02137_),
    .Y(_03892_));
 sky130_fd_sc_hd__o211ai_1 _21489_ (.A1(_02057_),
    .A2(_02183_),
    .B1(_03892_),
    .C1(net3745),
    .Y(_03893_));
 sky130_fd_sc_hd__a221oi_4 _21490_ (.A1(net3503),
    .A2(_02006_),
    .B1(net3603),
    .B2(_02221_),
    .C1(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__a21oi_2 _21491_ (.A1(net3756),
    .A2(_03888_),
    .B1(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_4 _21492_ (.A(net3738),
    .B(_11404_),
    .Y(_03896_));
 sky130_fd_sc_hd__o21ai_4 _21493_ (.A1(net3738),
    .A2(_03895_),
    .B1(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__mux4_2 _21494_ (.A0(net41),
    .A1(net55),
    .A2(\load_store_unit_i.rdata_q[22] ),
    .A3(net32),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03898_));
 sky130_fd_sc_hd__a21oi_1 _21495_ (.A1(_01670_),
    .A2(_03898_),
    .B1(_03289_),
    .Y(_03899_));
 sky130_fd_sc_hd__a21oi_2 _21496_ (.A1(net3469),
    .A2(_03897_),
    .B1(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_419 ();
 sky130_fd_sc_hd__mux2_1 _21498_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .A1(net3412),
    .S(_03095_),
    .X(_00529_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_418 ();
 sky130_fd_sc_hd__xor2_2 _21500_ (.A(net3531),
    .B(_02287_),
    .X(_03903_));
 sky130_fd_sc_hd__and2_4 _21501_ (.A(net3670),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__or2_0 _21502_ (.A(_03670_),
    .B(_03755_),
    .X(_03905_));
 sky130_fd_sc_hd__o21ai_0 _21503_ (.A1(net3465),
    .A2(_03668_),
    .B1(_03757_),
    .Y(_03906_));
 sky130_fd_sc_hd__a21boi_0 _21504_ (.A1(_03905_),
    .A2(_03906_),
    .B1_N(_03881_),
    .Y(_03907_));
 sky130_fd_sc_hd__inv_1 _21505_ (.A(_03872_),
    .Y(_03908_));
 sky130_fd_sc_hd__maj3_2 _21506_ (.A(_03876_),
    .B(_03908_),
    .C(_03877_),
    .X(_03909_));
 sky130_fd_sc_hd__nor2_1 _21507_ (.A(_03850_),
    .B(_03870_),
    .Y(_03910_));
 sky130_fd_sc_hd__nor2_1 _21508_ (.A(_03783_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__a21oi_2 _21509_ (.A1(_03850_),
    .A2(_03870_),
    .B1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__maj3_1 _21510_ (.A(_03828_),
    .B(_03813_),
    .C(_03829_),
    .X(_03913_));
 sky130_fd_sc_hd__inv_1 _21511_ (.A(_03856_),
    .Y(_03914_));
 sky130_fd_sc_hd__nor2_1 _21512_ (.A(_03914_),
    .B(_03867_),
    .Y(_03915_));
 sky130_fd_sc_hd__maj3_1 _21513_ (.A(_03858_),
    .B(_03859_),
    .C(_03860_),
    .X(_03916_));
 sky130_fd_sc_hd__nor2_1 _21514_ (.A(_02240_),
    .B(net3632),
    .Y(_03917_));
 sky130_fd_sc_hd__nor2_1 _21515_ (.A(net3639),
    .B(_02856_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor2_1 _21516_ (.A(_02243_),
    .B(_03188_),
    .Y(_03919_));
 sky130_fd_sc_hd__xor2_1 _21517_ (.A(_03918_),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__xor2_1 _21518_ (.A(_03917_),
    .B(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__maj3_1 _21519_ (.A(_03822_),
    .B(_03823_),
    .C(_03824_),
    .X(_03922_));
 sky130_fd_sc_hd__xor2_1 _21520_ (.A(_03921_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__xor2_1 _21521_ (.A(_03916_),
    .B(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__maj3_1 _21522_ (.A(_03863_),
    .B(_03862_),
    .C(_03865_),
    .X(_03925_));
 sky130_fd_sc_hd__xor2_1 _21523_ (.A(_03924_),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__xnor2_1 _21524_ (.A(_03915_),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__xnor2_1 _21525_ (.A(_03913_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__nor2_2 _21526_ (.A(net3636),
    .B(_02744_),
    .Y(_03929_));
 sky130_fd_sc_hd__nor2_1 _21527_ (.A(net3635),
    .B(net3633),
    .Y(_03930_));
 sky130_fd_sc_hd__nor2_1 _21528_ (.A(net3638),
    .B(_02877_),
    .Y(_03931_));
 sky130_fd_sc_hd__xor2_1 _21529_ (.A(_03930_),
    .B(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__xnor2_1 _21530_ (.A(_03929_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__maj3_1 _21531_ (.A(_03815_),
    .B(_03816_),
    .C(_03817_),
    .X(_03934_));
 sky130_fd_sc_hd__nor2_1 _21532_ (.A(_02505_),
    .B(net3634),
    .Y(_03935_));
 sky130_fd_sc_hd__nor2_1 _21533_ (.A(_02476_),
    .B(_02764_),
    .Y(_03936_));
 sky130_fd_sc_hd__nor2_1 _21534_ (.A(_02334_),
    .B(_02680_),
    .Y(_03937_));
 sky130_fd_sc_hd__xor2_1 _21535_ (.A(_03936_),
    .B(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__xnor2_1 _21536_ (.A(_03935_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__xor2_1 _21537_ (.A(_03934_),
    .B(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__xnor2_1 _21538_ (.A(_03933_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2b_2 _21539_ (.A(_03787_),
    .B_N(_03788_),
    .Y(_03942_));
 sky130_fd_sc_hd__o32ai_4 _21540_ (.A1(_03785_),
    .A2(_03786_),
    .A3(_03788_),
    .B1(_03942_),
    .B2(_03707_),
    .Y(_03943_));
 sky130_fd_sc_hd__maj3_1 _21541_ (.A(_03821_),
    .B(_03819_),
    .C(_03826_),
    .X(_03944_));
 sky130_fd_sc_hd__xor2_1 _21542_ (.A(_03943_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__xnor2_1 _21543_ (.A(_03941_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__nand3_2 _21544_ (.A(_01757_),
    .B(_01780_),
    .C(_03570_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _21545_ (.A(_01783_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__o21ai_2 _21546_ (.A1(_01757_),
    .A2(_01780_),
    .B1(net3646),
    .Y(_03949_));
 sky130_fd_sc_hd__a21oi_4 _21547_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_02987_),
    .Y(_03950_));
 sky130_fd_sc_hd__xnor2_4 _21548_ (.A(_03707_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__xnor2_4 _21549_ (.A(_03575_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__a21o_4 _21550_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(_03681_),
    .B1(_03471_),
    .X(_03953_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_417 ();
 sky130_fd_sc_hd__a21oi_2 _21552_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_03681_),
    .B1(_03471_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _21553_ (.A(_03460_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nor2_2 _21554_ (.A(_03460_),
    .B(_03955_),
    .Y(_03957_));
 sky130_fd_sc_hd__a21oi_2 _21555_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_10746_),
    .B1(_03310_),
    .Y(_03958_));
 sky130_fd_sc_hd__o21ai_0 _21556_ (.A1(_03685_),
    .A2(_03958_),
    .B1(_03460_),
    .Y(_03959_));
 sky130_fd_sc_hd__a221oi_1 _21557_ (.A1(_03792_),
    .A2(_03957_),
    .B1(_03959_),
    .B2(net3629),
    .C1(_03691_),
    .Y(_03960_));
 sky130_fd_sc_hd__a21oi_1 _21558_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_03681_),
    .B1(_03471_),
    .Y(_03961_));
 sky130_fd_sc_hd__nor2_1 _21559_ (.A(net3627),
    .B(_03796_),
    .Y(_03962_));
 sky130_fd_sc_hd__o21ai_0 _21560_ (.A1(_03792_),
    .A2(_03796_),
    .B1(net3627),
    .Y(_03963_));
 sky130_fd_sc_hd__a221oi_1 _21561_ (.A1(_03961_),
    .A2(_03962_),
    .B1(_03963_),
    .B2(_03459_),
    .C1(_03803_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand2_1 _21562_ (.A(net3629),
    .B(_03957_),
    .Y(_03965_));
 sky130_fd_sc_hd__o221ai_2 _21563_ (.A1(net3629),
    .A2(_03956_),
    .B1(_03960_),
    .B2(_03964_),
    .C1(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__xnor2_2 _21564_ (.A(_03953_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__xor2_1 _21565_ (.A(_03952_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__xnor2_1 _21566_ (.A(_03946_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__maj3_1 _21567_ (.A(_03791_),
    .B(_03798_),
    .C(_03810_),
    .X(_03970_));
 sky130_fd_sc_hd__xnor2_1 _21568_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__maj3_1 _21569_ (.A(_03811_),
    .B(_03831_),
    .C(_03848_),
    .X(_03972_));
 sky130_fd_sc_hd__xor2_1 _21570_ (.A(_03971_),
    .B(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__xnor2_1 _21571_ (.A(_03928_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _21572_ (.A(_03852_),
    .B(_03868_),
    .Y(_03975_));
 sky130_fd_sc_hd__nor2_1 _21573_ (.A(_03852_),
    .B(_03868_),
    .Y(_03976_));
 sky130_fd_sc_hd__a21oi_1 _21574_ (.A1(_03853_),
    .A2(_03975_),
    .B1(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__nor2_1 _21575_ (.A(_03974_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__and2_0 _21576_ (.A(_03974_),
    .B(_03977_),
    .X(_03979_));
 sky130_fd_sc_hd__nor2_1 _21577_ (.A(_03978_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__xor2_1 _21578_ (.A(_03912_),
    .B(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__xnor2_1 _21579_ (.A(_03909_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21ai_0 _21580_ (.A1(_03880_),
    .A2(_03907_),
    .B1(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__or3_1 _21581_ (.A(_03880_),
    .B(_03907_),
    .C(_03982_),
    .X(_03984_));
 sky130_fd_sc_hd__a21oi_2 _21582_ (.A1(_03983_),
    .A2(_03984_),
    .B1(net3670),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2b_2 _21583_ (.A_N(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B(net3937),
    .Y(_03986_));
 sky130_fd_sc_hd__o31ai_4 _21584_ (.A1(net3937),
    .A2(_03904_),
    .A3(_03985_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _21585_ (.A(_09907_),
    .B(_09937_),
    .Y(_03988_));
 sky130_fd_sc_hd__xor2_1 _21586_ (.A(_02133_),
    .B(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__o21ai_0 _21587_ (.A1(_09907_),
    .A2(_09937_),
    .B1(_02137_),
    .Y(_03990_));
 sky130_fd_sc_hd__a21oi_1 _21588_ (.A1(_02127_),
    .A2(_03989_),
    .B1(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a221oi_2 _21589_ (.A1(net3602),
    .A2(_02064_),
    .B1(_02121_),
    .B2(net3603),
    .C1(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__o21ai_4 _21590_ (.A1(net3504),
    .A2(_02702_),
    .B1(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__nor2_2 _21591_ (.A(net3756),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__a21oi_4 _21592_ (.A1(net3756),
    .A2(_03987_),
    .B1(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_2 _21593_ (.A(_11423_),
    .B(net3469),
    .Y(_03996_));
 sky130_fd_sc_hd__mux4_2 _21594_ (.A0(net42),
    .A1(net56),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .A3(net33),
    .S0(net3822),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03997_));
 sky130_fd_sc_hd__a21o_1 _21595_ (.A1(_01670_),
    .A2(_03997_),
    .B1(_03289_),
    .X(_03998_));
 sky130_fd_sc_hd__o21ai_2 _21596_ (.A1(_03995_),
    .A2(_03996_),
    .B1(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_416 ();
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .B(_02153_),
    .Y(_04001_));
 sky130_fd_sc_hd__o21ai_0 _21599_ (.A1(_02153_),
    .A2(net3411),
    .B1(_04001_),
    .Y(_00530_));
 sky130_fd_sc_hd__nor2_1 _21600_ (.A(_02423_),
    .B(_01662_),
    .Y(_04002_));
 sky130_fd_sc_hd__a211oi_2 _21601_ (.A1(_02423_),
    .A2(_01664_),
    .B1(_02847_),
    .C1(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _21602_ (.A(net3670),
    .B(_01998_),
    .Y(_04004_));
 sky130_fd_sc_hd__inv_1 _21603_ (.A(_03909_),
    .Y(_04005_));
 sky130_fd_sc_hd__nor2_1 _21604_ (.A(_03756_),
    .B(_03880_),
    .Y(_04006_));
 sky130_fd_sc_hd__o21ai_1 _21605_ (.A1(_04005_),
    .A2(_03981_),
    .B1(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_1 _21606_ (.A(net3488),
    .B(_03515_),
    .Y(_04008_));
 sky130_fd_sc_hd__a21o_1 _21607_ (.A1(_03395_),
    .A2(_04008_),
    .B1(_03538_),
    .X(_04009_));
 sky130_fd_sc_hd__o311ai_1 _21608_ (.A1(_03299_),
    .A2(_03419_),
    .A3(_03538_),
    .B1(_03637_),
    .C1(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__a21oi_1 _21609_ (.A1(_03638_),
    .A2(net3467),
    .B1(_03758_),
    .Y(_04011_));
 sky130_fd_sc_hd__xnor2_1 _21610_ (.A(_03912_),
    .B(_03980_),
    .Y(_04012_));
 sky130_fd_sc_hd__maj3_1 _21611_ (.A(_03881_),
    .B(_03909_),
    .C(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__o21ai_0 _21612_ (.A1(_04007_),
    .A2(_04011_),
    .B1(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__o21bai_1 _21613_ (.A1(_03912_),
    .A2(_03979_),
    .B1_N(_03978_),
    .Y(_04015_));
 sky130_fd_sc_hd__maj3_1 _21614_ (.A(_03915_),
    .B(_03913_),
    .C(_03926_),
    .X(_04016_));
 sky130_fd_sc_hd__inv_1 _21615_ (.A(_03972_),
    .Y(_04017_));
 sky130_fd_sc_hd__maj3_1 _21616_ (.A(_03928_),
    .B(_03971_),
    .C(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__maj3_1 _21617_ (.A(_03941_),
    .B(_03943_),
    .C(_03944_),
    .X(_04019_));
 sky130_fd_sc_hd__nor2_2 _21618_ (.A(_03924_),
    .B(_03925_),
    .Y(_04020_));
 sky130_fd_sc_hd__nor2_1 _21619_ (.A(_02334_),
    .B(_02784_),
    .Y(_04021_));
 sky130_fd_sc_hd__nor2_1 _21620_ (.A(_02240_),
    .B(_02856_),
    .Y(_04022_));
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(net3637),
    .B(_03060_),
    .Y(_04023_));
 sky130_fd_sc_hd__xor2_1 _21622_ (.A(_04022_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__xor2_1 _21623_ (.A(_04021_),
    .B(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__maj3_1 _21624_ (.A(_03917_),
    .B(_03918_),
    .C(_03919_),
    .X(_04026_));
 sky130_fd_sc_hd__maj3_1 _21625_ (.A(_03936_),
    .B(_03935_),
    .C(_03937_),
    .X(_04027_));
 sky130_fd_sc_hd__xnor2_1 _21626_ (.A(_04026_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_1 _21627_ (.A(_04025_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _21628_ (.A(_03921_),
    .B(_03922_),
    .Y(_04030_));
 sky130_fd_sc_hd__nor2_1 _21629_ (.A(_03921_),
    .B(_03922_),
    .Y(_04031_));
 sky130_fd_sc_hd__a21oi_2 _21630_ (.A1(_03916_),
    .A2(_04030_),
    .B1(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__xnor2_1 _21631_ (.A(_04029_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__xor2_1 _21632_ (.A(_04020_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__xnor2_1 _21633_ (.A(_04019_),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__inv_1 _21634_ (.A(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_415 ();
 sky130_fd_sc_hd__inv_6 _21636_ (.A(_03575_),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_2 _21637_ (.A(_04038_),
    .B(_03951_),
    .Y(_04039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_414 ();
 sky130_fd_sc_hd__a21oi_1 _21639_ (.A1(net3627),
    .A2(_03958_),
    .B1(net3629),
    .Y(_04041_));
 sky130_fd_sc_hd__a21oi_2 _21640_ (.A1(_03460_),
    .A2(_03796_),
    .B1(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__a21oi_1 _21641_ (.A1(_03792_),
    .A2(_03962_),
    .B1(_03957_),
    .Y(_04043_));
 sky130_fd_sc_hd__o32ai_1 _21642_ (.A1(_03470_),
    .A2(_03961_),
    .A3(_03796_),
    .B1(_04043_),
    .B2(_03459_),
    .Y(_04044_));
 sky130_fd_sc_hd__a21oi_1 _21643_ (.A1(net3627),
    .A2(_03685_),
    .B1(net3629),
    .Y(_04045_));
 sky130_fd_sc_hd__a21oi_1 _21644_ (.A1(_03460_),
    .A2(_03792_),
    .B1(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor3_1 _21645_ (.A(_03691_),
    .B(_03955_),
    .C(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__a21oi_1 _21646_ (.A1(_03691_),
    .A2(_04044_),
    .B1(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_1 _21647_ (.A(_03953_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__a31oi_2 _21648_ (.A1(_03803_),
    .A2(_03953_),
    .A3(_04042_),
    .B1(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__xnor2_4 _21649_ (.A(_03564_),
    .B(_03950_),
    .Y(_04051_));
 sky130_fd_sc_hd__xnor2_1 _21650_ (.A(_04051_),
    .B(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_413 ();
 sky130_fd_sc_hd__nor2_1 _21652_ (.A(_03951_),
    .B(_03967_),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2_1 _21653_ (.A(_04050_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__o221a_1 _21654_ (.A1(_04039_),
    .A2(_04050_),
    .B1(_04052_),
    .B2(_04038_),
    .C1(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__maj3_1 _21655_ (.A(_03930_),
    .B(_03929_),
    .C(_03931_),
    .X(_04057_));
 sky130_fd_sc_hd__nand2b_2 _21656_ (.A_N(_02744_),
    .B(_02320_),
    .Y(_04058_));
 sky130_fd_sc_hd__nor2_1 _21657_ (.A(net3638),
    .B(_02987_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand2_1 _21658_ (.A(_02270_),
    .B(_03570_),
    .Y(_04060_));
 sky130_fd_sc_hd__xnor2_1 _21659_ (.A(_04059_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__xnor2_1 _21660_ (.A(_04058_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__nor2_1 _21661_ (.A(_02764_),
    .B(net3634),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2b_1 _21662_ (.A_N(_02476_),
    .B(_02900_),
    .Y(_04064_));
 sky130_fd_sc_hd__or2_4 _21663_ (.A(_02505_),
    .B(net3633),
    .X(_04065_));
 sky130_fd_sc_hd__xnor2_1 _21664_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__xnor2_1 _21665_ (.A(_04063_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__xnor3_1 _21666_ (.A(_04057_),
    .B(_04062_),
    .C(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__a21oi_2 _21667_ (.A1(_03564_),
    .A2(_03947_),
    .B1(net3646),
    .Y(_04069_));
 sky130_fd_sc_hd__a21oi_1 _21668_ (.A1(net3643),
    .A2(net3647),
    .B1(_03564_),
    .Y(_04070_));
 sky130_fd_sc_hd__o21ai_4 _21669_ (.A1(_04069_),
    .A2(_04070_),
    .B1(net3630),
    .Y(_04071_));
 sky130_fd_sc_hd__clkinvlp_4 _21670_ (.A(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _21671_ (.A(_03933_),
    .B(_03939_),
    .Y(_04073_));
 sky130_fd_sc_hd__nor2_1 _21672_ (.A(_03933_),
    .B(_03939_),
    .Y(_04074_));
 sky130_fd_sc_hd__a21oi_1 _21673_ (.A1(_03934_),
    .A2(_04073_),
    .B1(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__xnor2_1 _21674_ (.A(_04072_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__xnor2_2 _21675_ (.A(_04068_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__a21oi_4 _21676_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(_10746_),
    .B1(net3669),
    .Y(_04078_));
 sky130_fd_sc_hd__a21oi_2 _21677_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(_10746_),
    .B1(_03310_),
    .Y(_04079_));
 sky130_fd_sc_hd__o21ai_0 _21678_ (.A1(_03958_),
    .A2(_04079_),
    .B1(_03460_),
    .Y(_04080_));
 sky130_fd_sc_hd__a22o_1 _21679_ (.A1(_03953_),
    .A2(_03957_),
    .B1(_04080_),
    .B2(net3629),
    .X(_04081_));
 sky130_fd_sc_hd__nand2_1 _21680_ (.A(_03803_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__a21oi_1 _21681_ (.A1(_03958_),
    .A2(_04079_),
    .B1(_03460_),
    .Y(_04083_));
 sky130_fd_sc_hd__o22ai_1 _21682_ (.A1(_03953_),
    .A2(_03956_),
    .B1(_04083_),
    .B2(net3629),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _21683_ (.A(_03691_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__a21o_4 _21684_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(_10746_),
    .B1(net3669),
    .X(_04086_));
 sky130_fd_sc_hd__nand3_1 _21685_ (.A(net3629),
    .B(net3627),
    .C(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand3_1 _21686_ (.A(_03459_),
    .B(_03460_),
    .C(_04079_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand4_1 _21687_ (.A(_04082_),
    .B(_04085_),
    .C(_04087_),
    .D(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__xnor2_1 _21688_ (.A(_04078_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__xnor2_1 _21689_ (.A(_04077_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__xnor2_1 _21690_ (.A(_04056_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__xnor2_1 _21691_ (.A(_04036_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__maj3_1 _21692_ (.A(_03946_),
    .B(_03968_),
    .C(_03970_),
    .X(_04094_));
 sky130_fd_sc_hd__xnor2_1 _21693_ (.A(_04093_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__xnor3_1 _21694_ (.A(_04016_),
    .B(_04018_),
    .C(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_2 _21695_ (.A(_04015_),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__nor2_1 _21696_ (.A(_04015_),
    .B(_04096_),
    .Y(_04098_));
 sky130_fd_sc_hd__inv_1 _21697_ (.A(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _21698_ (.A(_04097_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__xnor2_1 _21699_ (.A(_04014_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_2 _21700_ (.A(_02000_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_4 _21701_ (.A(_04004_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__mux2i_4 _21702_ (.A0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A1(_04103_),
    .S(_08009_),
    .Y(_04104_));
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(net3557),
    .B(_02079_),
    .Y(_04105_));
 sky130_fd_sc_hd__nor2_4 _21704_ (.A(_02182_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__mux2i_2 _21705_ (.A0(_02108_),
    .A1(_03263_),
    .S(net3621),
    .Y(_04107_));
 sky130_fd_sc_hd__mux2i_1 _21706_ (.A0(_04107_),
    .A1(_02204_),
    .S(net3578),
    .Y(_04108_));
 sky130_fd_sc_hd__mux2i_1 _21707_ (.A0(_02449_),
    .A1(_04108_),
    .S(net3558),
    .Y(_04109_));
 sky130_fd_sc_hd__nor2_1 _21708_ (.A(_02056_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__a211oi_1 _21709_ (.A1(_02056_),
    .A2(_02949_),
    .B1(_04110_),
    .C1(net3557),
    .Y(_04111_));
 sky130_fd_sc_hd__o21bai_4 _21710_ (.A1(net3560),
    .A2(_02061_),
    .B1_N(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _21711_ (.A(_09987_),
    .B(_10018_),
    .Y(_04113_));
 sky130_fd_sc_hd__xor2_1 _21712_ (.A(_02133_),
    .B(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__a21oi_1 _21713_ (.A1(_09987_),
    .A2(_10018_),
    .B1(_03273_),
    .Y(_04115_));
 sky130_fd_sc_hd__o21ai_0 _21714_ (.A1(_02184_),
    .A2(_04114_),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand3_1 _21715_ (.A(net3746),
    .B(_08501_),
    .C(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__a21oi_1 _21716_ (.A1(net3603),
    .A2(_04112_),
    .B1(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__o21ai_2 _21717_ (.A1(_02057_),
    .A2(_04106_),
    .B1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a21oi_4 _21718_ (.A1(net273),
    .A2(_02006_),
    .B1(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__a221oi_1 _21719_ (.A1(net3738),
    .A2(_11439_),
    .B1(_04104_),
    .B2(net3756),
    .C1(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__o22ai_2 _21720_ (.A1(_03289_),
    .A2(_04003_),
    .B1(_04121_),
    .B2(net3472),
    .Y(_04122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_412 ();
 sky130_fd_sc_hd__nand2_1 _21722_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .B(_02153_),
    .Y(_04124_));
 sky130_fd_sc_hd__o21ai_0 _21723_ (.A1(_02153_),
    .A2(net3410),
    .B1(_04124_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand3_1 _21724_ (.A(_03757_),
    .B(_03881_),
    .C(_04005_),
    .Y(_04125_));
 sky130_fd_sc_hd__a221o_1 _21725_ (.A1(_03756_),
    .A2(_03881_),
    .B1(_04012_),
    .B2(_04125_),
    .C1(_03880_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_1 _21726_ (.A1(_03757_),
    .A2(_03881_),
    .B1(_03880_),
    .Y(_04127_));
 sky130_fd_sc_hd__maj3_1 _21727_ (.A(_04005_),
    .B(_03981_),
    .C(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__nor2_1 _21728_ (.A(_04098_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__o31ai_2 _21729_ (.A1(_03666_),
    .A2(_03668_),
    .A3(_04126_),
    .B1(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _21730_ (.A(_04097_),
    .B(net3458),
    .Y(_04131_));
 sky130_fd_sc_hd__maj3_2 _21731_ (.A(_04016_),
    .B(_04018_),
    .C(_04095_),
    .X(_04132_));
 sky130_fd_sc_hd__nand2_1 _21732_ (.A(_04019_),
    .B(_04033_),
    .Y(_04133_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_04019_),
    .B(_04033_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21oi_1 _21734_ (.A1(_04020_),
    .A2(_04133_),
    .B1(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__inv_1 _21735_ (.A(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__nor3_1 _21736_ (.A(net3627),
    .B(_03958_),
    .C(_04086_),
    .Y(_04137_));
 sky130_fd_sc_hd__a21oi_1 _21737_ (.A1(net3627),
    .A2(_04086_),
    .B1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__o32ai_1 _21738_ (.A1(_03470_),
    .A2(_03958_),
    .A3(_04086_),
    .B1(_04138_),
    .B2(_03459_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand3_1 _21739_ (.A(_03691_),
    .B(_04078_),
    .C(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__o21ai_0 _21740_ (.A1(_03460_),
    .A2(_04086_),
    .B1(_03459_),
    .Y(_04141_));
 sky130_fd_sc_hd__o21ai_1 _21741_ (.A1(net3627),
    .A2(_04079_),
    .B1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand2_1 _21742_ (.A(_04086_),
    .B(_04078_),
    .Y(_04143_));
 sky130_fd_sc_hd__o22ai_1 _21743_ (.A1(_04078_),
    .A2(_04142_),
    .B1(_04143_),
    .B2(_04042_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _21744_ (.A(_03803_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_4 _21745_ (.A(_04140_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__xnor2_1 _21746_ (.A(_04051_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nor2_1 _21747_ (.A(_04038_),
    .B(_04051_),
    .Y(_04148_));
 sky130_fd_sc_hd__nor3_1 _21748_ (.A(_03951_),
    .B(_04090_),
    .C(_04146_),
    .Y(_04149_));
 sky130_fd_sc_hd__a221oi_1 _21749_ (.A1(_04038_),
    .A2(_04147_),
    .B1(_04148_),
    .B2(_04146_),
    .C1(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21oi_1 _21750_ (.A1(_02503_),
    .A2(_02744_),
    .B1(_02270_),
    .Y(_04151_));
 sky130_fd_sc_hd__a21oi_1 _21751_ (.A1(_02744_),
    .A2(_02987_),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__or3_4 _21752_ (.A(net3635),
    .B(_02877_),
    .C(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _21753_ (.A(net3638),
    .B(net3636),
    .Y(_04154_));
 sky130_fd_sc_hd__nand3_1 _21754_ (.A(_02320_),
    .B(_02744_),
    .C(_03570_),
    .Y(_04155_));
 sky130_fd_sc_hd__o2111ai_1 _21755_ (.A1(net3638),
    .A2(_04058_),
    .B1(_04154_),
    .C1(_04155_),
    .D1(net3630),
    .Y(_04156_));
 sky130_fd_sc_hd__nor2_1 _21756_ (.A(net3634),
    .B(_02680_),
    .Y(_04157_));
 sky130_fd_sc_hd__nor2_1 _21757_ (.A(_02764_),
    .B(net3633),
    .Y(_04158_));
 sky130_fd_sc_hd__nor2_1 _21758_ (.A(_02505_),
    .B(_02744_),
    .Y(_04159_));
 sky130_fd_sc_hd__xor2_1 _21759_ (.A(_04158_),
    .B(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__xnor2_1 _21760_ (.A(_04157_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__a21oi_2 _21761_ (.A1(_04153_),
    .A2(_04156_),
    .B1(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__and3_1 _21762_ (.A(_04153_),
    .B(_04156_),
    .C(_04161_),
    .X(_04163_));
 sky130_fd_sc_hd__nor2_2 _21763_ (.A(_04162_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__maj3_1 _21764_ (.A(_04057_),
    .B(_04062_),
    .C(_04067_),
    .X(_04165_));
 sky130_fd_sc_hd__xor2_1 _21765_ (.A(_04071_),
    .B(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__xnor2_2 _21766_ (.A(_04164_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_411 ();
 sky130_fd_sc_hd__a21oi_4 _21768_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(_03681_),
    .B1(net3731),
    .Y(_04169_));
 sky130_fd_sc_hd__a21oi_2 _21769_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(_03681_),
    .B1(net3731),
    .Y(_04170_));
 sky130_fd_sc_hd__nor3_1 _21770_ (.A(_03459_),
    .B(_03460_),
    .C(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__a21o_4 _21771_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(_03681_),
    .B1(_03471_),
    .X(_04172_));
 sky130_fd_sc_hd__nor3_1 _21772_ (.A(net3629),
    .B(net3627),
    .C(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__nand2_1 _21773_ (.A(_03953_),
    .B(_04172_),
    .Y(_04174_));
 sky130_fd_sc_hd__maj3_1 _21774_ (.A(_03459_),
    .B(_03460_),
    .C(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__o21ai_0 _21775_ (.A1(_03953_),
    .A2(_04172_),
    .B1(net3627),
    .Y(_04176_));
 sky130_fd_sc_hd__nor3_1 _21776_ (.A(net3627),
    .B(_03953_),
    .C(_04172_),
    .Y(_04177_));
 sky130_fd_sc_hd__a21oi_1 _21777_ (.A1(_03459_),
    .A2(_04176_),
    .B1(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__mux2i_1 _21778_ (.A0(_04175_),
    .A1(_04178_),
    .S(_03691_),
    .Y(_04179_));
 sky130_fd_sc_hd__nor3_2 _21779_ (.A(_04171_),
    .B(_04173_),
    .C(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__xnor2_2 _21780_ (.A(_04169_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__xnor2_1 _21781_ (.A(_04167_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__xnor2_1 _21782_ (.A(_04150_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_2 _21783_ (.A(_04029_),
    .B(_04032_),
    .Y(_04184_));
 sky130_fd_sc_hd__maj3_1 _21784_ (.A(_04071_),
    .B(_04068_),
    .C(_04075_),
    .X(_04185_));
 sky130_fd_sc_hd__nor2_1 _21785_ (.A(_02476_),
    .B(_02784_),
    .Y(_04186_));
 sky130_fd_sc_hd__nor2_1 _21786_ (.A(_02334_),
    .B(_02856_),
    .Y(_04187_));
 sky130_fd_sc_hd__nor2b_2 _21787_ (.A(_03188_),
    .B_N(_02240_),
    .Y(_04188_));
 sky130_fd_sc_hd__xnor2_1 _21788_ (.A(_04187_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__xnor2_1 _21789_ (.A(_04186_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__maj3_1 _21790_ (.A(_04021_),
    .B(_04022_),
    .C(_04023_),
    .X(_04191_));
 sky130_fd_sc_hd__inv_1 _21791_ (.A(_04064_),
    .Y(_04192_));
 sky130_fd_sc_hd__inv_1 _21792_ (.A(_04065_),
    .Y(_04193_));
 sky130_fd_sc_hd__maj3_1 _21793_ (.A(_04192_),
    .B(_04063_),
    .C(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__xnor2_1 _21794_ (.A(_04191_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__xnor2_1 _21795_ (.A(_04190_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__maj3_2 _21796_ (.A(_04026_),
    .B(_04025_),
    .C(_04027_),
    .X(_04197_));
 sky130_fd_sc_hd__xnor2_1 _21797_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__xnor2_1 _21798_ (.A(_04185_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__xor2_1 _21799_ (.A(_04184_),
    .B(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__xor2_1 _21800_ (.A(_04183_),
    .B(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_410 ();
 sky130_fd_sc_hd__nand2_1 _21802_ (.A(_04051_),
    .B(_04090_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _21803_ (.A(_04077_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand3_1 _21804_ (.A(net3629),
    .B(net3627),
    .C(_03953_),
    .Y(_04205_));
 sky130_fd_sc_hd__or3_1 _21805_ (.A(net3629),
    .B(net3627),
    .C(_03953_),
    .X(_04206_));
 sky130_fd_sc_hd__mux2i_1 _21806_ (.A0(_04081_),
    .A1(_04084_),
    .S(_03691_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand3_1 _21807_ (.A(_04205_),
    .B(_04206_),
    .C(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__xnor2_1 _21808_ (.A(_04170_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__nor2_1 _21809_ (.A(_04051_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__a211oi_1 _21810_ (.A1(_03967_),
    .A2(_04204_),
    .B1(_04210_),
    .C1(_04038_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2b_1 _21811_ (.A_N(_04209_),
    .B(_04051_),
    .Y(_04212_));
 sky130_fd_sc_hd__a21oi_1 _21812_ (.A1(_04077_),
    .A2(_04212_),
    .B1(_03967_),
    .Y(_04213_));
 sky130_fd_sc_hd__a211oi_1 _21813_ (.A1(_03951_),
    .A2(_04209_),
    .B1(_04213_),
    .C1(net3571),
    .Y(_04214_));
 sky130_fd_sc_hd__o22ai_1 _21814_ (.A1(_04051_),
    .A2(_04077_),
    .B1(_04211_),
    .B2(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__xnor2_1 _21815_ (.A(_03952_),
    .B(_04209_),
    .Y(_04216_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_04077_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__a21oi_2 _21817_ (.A1(_04050_),
    .A2(_04215_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__xor2_1 _21818_ (.A(_04201_),
    .B(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__maj3_1 _21819_ (.A(_04036_),
    .B(_04092_),
    .C(_04094_),
    .X(_04220_));
 sky130_fd_sc_hd__xnor3_1 _21820_ (.A(_04136_),
    .B(_04219_),
    .C(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__xnor2_1 _21821_ (.A(_04132_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__xnor2_1 _21822_ (.A(_04131_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2_2 _21823_ (.A(_02000_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__o21ai_4 _21824_ (.A1(_02000_),
    .A2(_02289_),
    .B1(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__mux2i_1 _21825_ (.A0(_03264_),
    .A1(_02111_),
    .S(net3578),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _21826_ (.A(net3558),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__o21ai_0 _21827_ (.A1(net3558),
    .A2(_02393_),
    .B1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _21828_ (.A(_02016_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__o211ai_1 _21829_ (.A1(_02016_),
    .A2(_02824_),
    .B1(_04229_),
    .C1(net3560),
    .Y(_04230_));
 sky130_fd_sc_hd__o21ai_2 _21830_ (.A1(net3560),
    .A2(_02180_),
    .B1(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__nor2_2 _21831_ (.A(net3557),
    .B(_02219_),
    .Y(_04232_));
 sky130_fd_sc_hd__nor2_2 _21832_ (.A(_02063_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__a22oi_2 _21833_ (.A1(net3603),
    .A2(_04231_),
    .B1(_04233_),
    .B2(net3602),
    .Y(_04234_));
 sky130_fd_sc_hd__nor2_1 _21834_ (.A(_10060_),
    .B(_10098_),
    .Y(_04235_));
 sky130_fd_sc_hd__xor2_1 _21835_ (.A(_02133_),
    .B(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__a21oi_1 _21836_ (.A1(_10060_),
    .A2(_10098_),
    .B1(_03273_),
    .Y(_04237_));
 sky130_fd_sc_hd__o21ai_2 _21837_ (.A1(_02184_),
    .A2(_04236_),
    .B1(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand3_4 _21838_ (.A(net3737),
    .B(_04234_),
    .C(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__a21oi_1 _21839_ (.A1(net3495),
    .A2(_02006_),
    .B1(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__nor2_1 _21840_ (.A(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .B(_13047_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_04240_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__o31ai_2 _21842_ (.A1(net3937),
    .A2(net3747),
    .A3(_04225_),
    .B1(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _21843_ (.A(net3822),
    .B(_02163_),
    .Y(_04244_));
 sky130_fd_sc_hd__o21ai_2 _21844_ (.A1(net3822),
    .A2(_02162_),
    .B1(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__a21oi_2 _21845_ (.A1(_01670_),
    .A2(_04245_),
    .B1(_03289_),
    .Y(_04246_));
 sky130_fd_sc_hd__a31o_4 _21846_ (.A1(_11455_),
    .A2(net3469),
    .A3(_04243_),
    .B1(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_409 ();
 sky130_fd_sc_hd__nand2_1 _21848_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .B(_02153_),
    .Y(_04249_));
 sky130_fd_sc_hd__o21ai_0 _21849_ (.A1(_02153_),
    .A2(net3409),
    .B1(_04249_),
    .Y(_00532_));
 sky130_fd_sc_hd__nor2_1 _21850_ (.A(_02000_),
    .B(_02383_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2b_2 _21851_ (.A_N(_04221_),
    .B(_04132_),
    .Y(_04251_));
 sky130_fd_sc_hd__o211ai_1 _21852_ (.A1(_04007_),
    .A2(_04011_),
    .B1(_04099_),
    .C1(_04013_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _21853_ (.A(_04097_),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2b_2 _21854_ (.A_N(_04132_),
    .B(_04221_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21boi_0 _21855_ (.A1(_04251_),
    .A2(_04253_),
    .B1_N(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__maj3_1 _21856_ (.A(_04136_),
    .B(_04219_),
    .C(_04220_),
    .X(_04256_));
 sky130_fd_sc_hd__maj3_1 _21857_ (.A(_04183_),
    .B(_04200_),
    .C(_04218_),
    .X(_04257_));
 sky130_fd_sc_hd__maj3_2 _21858_ (.A(_04184_),
    .B(_04185_),
    .C(_04198_),
    .X(_04258_));
 sky130_fd_sc_hd__xnor2_1 _21859_ (.A(_04038_),
    .B(_04181_),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _21860_ (.A(_03953_),
    .B(_04170_),
    .Y(_04260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_408 ();
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(net3627),
    .B(_04260_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21oi_1 _21863_ (.A1(net3627),
    .A2(_04172_),
    .B1(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o22ai_1 _21864_ (.A1(_03470_),
    .A2(_04260_),
    .B1(_04263_),
    .B2(_03459_),
    .Y(_04264_));
 sky130_fd_sc_hd__a21o_4 _21865_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(_03681_),
    .B1(net3731),
    .X(_04265_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_04170_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__o21ai_0 _21867_ (.A1(net3627),
    .A2(_04078_),
    .B1(net3629),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(net3627),
    .B(_04078_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21oi_4 _21869_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(_10746_),
    .B1(net3669),
    .Y(_04269_));
 sky130_fd_sc_hd__a21oi_1 _21870_ (.A1(_04267_),
    .A2(_04268_),
    .B1(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__a21oi_1 _21871_ (.A1(_04142_),
    .A2(_04266_),
    .B1(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__nor2_1 _21872_ (.A(net3577),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a31o_1 _21873_ (.A1(net3577),
    .A2(_04169_),
    .A3(_04264_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a21oi_2 _21874_ (.A1(_04051_),
    .A2(_04259_),
    .B1(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__o21ai_0 _21875_ (.A1(_02744_),
    .A2(_03570_),
    .B1(_04060_),
    .Y(_04275_));
 sky130_fd_sc_hd__a32o_1 _21876_ (.A1(_03570_),
    .A2(_02987_),
    .A3(_03929_),
    .B1(_04059_),
    .B2(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__a21oi_2 _21877_ (.A1(_02320_),
    .A2(_04276_),
    .B1(_04162_),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _21878_ (.A(_02764_),
    .B(_02744_),
    .Y(_04278_));
 sky130_fd_sc_hd__nor2_1 _21879_ (.A(_02505_),
    .B(_02877_),
    .Y(_04279_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(net3633),
    .B(_02680_),
    .Y(_04280_));
 sky130_fd_sc_hd__xor2_1 _21881_ (.A(_04279_),
    .B(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__xnor2_1 _21882_ (.A(_04278_),
    .B(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__xnor2_1 _21883_ (.A(_04277_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__o21ai_0 _21884_ (.A1(_02270_),
    .A2(_02877_),
    .B1(_02503_),
    .Y(_04284_));
 sky130_fd_sc_hd__o21ai_1 _21885_ (.A1(net3636),
    .A2(_03570_),
    .B1(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__nor2_2 _21886_ (.A(_02270_),
    .B(_02320_),
    .Y(_04286_));
 sky130_fd_sc_hd__a221o_4 _21887_ (.A1(_02320_),
    .A2(_04285_),
    .B1(_04286_),
    .B2(net3638),
    .C1(_02987_),
    .X(_04287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_407 ();
 sky130_fd_sc_hd__xor2_2 _21889_ (.A(_04071_),
    .B(_04287_),
    .X(_04289_));
 sky130_fd_sc_hd__xnor2_1 _21890_ (.A(_03952_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_1 _21891_ (.A(_04283_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__nor3_1 _21892_ (.A(net3627),
    .B(_04172_),
    .C(_04169_),
    .Y(_04292_));
 sky130_fd_sc_hd__a311oi_1 _21893_ (.A1(net3627),
    .A2(net3577),
    .A3(_04169_),
    .B1(_04292_),
    .C1(_03459_),
    .Y(_04293_));
 sky130_fd_sc_hd__nor3_1 _21894_ (.A(_03460_),
    .B(_04172_),
    .C(_04269_),
    .Y(_04294_));
 sky130_fd_sc_hd__a211oi_1 _21895_ (.A1(_03460_),
    .A2(_04169_),
    .B1(_04294_),
    .C1(net3629),
    .Y(_04295_));
 sky130_fd_sc_hd__o22ai_2 _21896_ (.A1(_03800_),
    .A2(_04266_),
    .B1(_04293_),
    .B2(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21oi_1 _21897_ (.A1(net3627),
    .A2(_04265_),
    .B1(net3629),
    .Y(_04297_));
 sky130_fd_sc_hd__a21oi_1 _21898_ (.A1(_03460_),
    .A2(_04269_),
    .B1(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__a21oi_4 _21899_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_10746_),
    .B1(net3669),
    .Y(_04299_));
 sky130_fd_sc_hd__xnor2_1 _21900_ (.A(_04298_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__xnor2_1 _21901_ (.A(_04296_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__xnor2_1 _21902_ (.A(_04291_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__xnor2_1 _21903_ (.A(_04274_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__nand2_2 _21904_ (.A(_04196_),
    .B(_04197_),
    .Y(_04304_));
 sky130_fd_sc_hd__maj3_1 _21905_ (.A(_04072_),
    .B(_04164_),
    .C(_04165_),
    .X(_04305_));
 sky130_fd_sc_hd__nor2_1 _21906_ (.A(net3634),
    .B(_02784_),
    .Y(_04306_));
 sky130_fd_sc_hd__nor2_1 _21907_ (.A(_02476_),
    .B(_02856_),
    .Y(_04307_));
 sky130_fd_sc_hd__nor2_2 _21908_ (.A(_03141_),
    .B(_03188_),
    .Y(_04308_));
 sky130_fd_sc_hd__xnor2_1 _21909_ (.A(_04307_),
    .B(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__xnor2_1 _21910_ (.A(_04306_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__maj3_1 _21911_ (.A(_04186_),
    .B(_04187_),
    .C(_04188_),
    .X(_04311_));
 sky130_fd_sc_hd__maj3_2 _21912_ (.A(_04158_),
    .B(_04157_),
    .C(_04159_),
    .X(_04312_));
 sky130_fd_sc_hd__xnor2_1 _21913_ (.A(_04311_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__xnor2_1 _21914_ (.A(_04310_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__maj3_1 _21915_ (.A(_04191_),
    .B(_04190_),
    .C(_04194_),
    .X(_04315_));
 sky130_fd_sc_hd__xor2_1 _21916_ (.A(_04314_),
    .B(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__nor2_1 _21917_ (.A(_04305_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_1 _21918_ (.A(_04305_),
    .B(_04316_),
    .Y(_04318_));
 sky130_fd_sc_hd__nor2b_1 _21919_ (.A(_04317_),
    .B_N(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__xnor2_1 _21920_ (.A(_04304_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__xor2_1 _21921_ (.A(_04303_),
    .B(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__xor2_1 _21922_ (.A(_03952_),
    .B(_04181_),
    .X(_04322_));
 sky130_fd_sc_hd__nor2_1 _21923_ (.A(_04167_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__nor3_1 _21924_ (.A(_04038_),
    .B(_04209_),
    .C(_04181_),
    .Y(_04324_));
 sky130_fd_sc_hd__and3_1 _21925_ (.A(_04038_),
    .B(_04209_),
    .C(_04181_),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _21926_ (.A(_03951_),
    .B(_04167_),
    .Y(_04326_));
 sky130_fd_sc_hd__o31ai_1 _21927_ (.A1(_03951_),
    .A2(_04324_),
    .A3(_04325_),
    .B1(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__nor2b_1 _21928_ (.A(_04167_),
    .B_N(_04090_),
    .Y(_04328_));
 sky130_fd_sc_hd__and3_1 _21929_ (.A(_03459_),
    .B(_03460_),
    .C(_04078_),
    .X(_04329_));
 sky130_fd_sc_hd__nor3_1 _21930_ (.A(_03459_),
    .B(_03460_),
    .C(_04078_),
    .Y(_04330_));
 sky130_fd_sc_hd__nor2_1 _21931_ (.A(_03691_),
    .B(_04175_),
    .Y(_04331_));
 sky130_fd_sc_hd__nor2_1 _21932_ (.A(_03803_),
    .B(_04178_),
    .Y(_04332_));
 sky130_fd_sc_hd__nor4_1 _21933_ (.A(_04329_),
    .B(_04330_),
    .C(_04331_),
    .D(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__xnor2_1 _21934_ (.A(_04269_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__nor2_1 _21935_ (.A(_04051_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21ai_0 _21936_ (.A1(_04328_),
    .A2(_04335_),
    .B1(_04038_),
    .Y(_04336_));
 sky130_fd_sc_hd__a2bb2o_1 _21937_ (.A1_N(_04090_),
    .A2_N(_04167_),
    .B1(_04334_),
    .B2(_03951_),
    .X(_04337_));
 sky130_fd_sc_hd__nand2_1 _21938_ (.A(net3571),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a31oi_1 _21939_ (.A1(_04327_),
    .A2(_04336_),
    .A3(_04338_),
    .B1(_04146_),
    .Y(_04339_));
 sky130_fd_sc_hd__nor2_2 _21940_ (.A(_04323_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__xnor2_1 _21941_ (.A(_04321_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__xnor2_1 _21942_ (.A(_04258_),
    .B(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__xnor2_1 _21943_ (.A(_04257_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__nand2_2 _21944_ (.A(_04256_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__or2_4 _21945_ (.A(_04256_),
    .B(_04343_),
    .X(_04345_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_406 ();
 sky130_fd_sc_hd__nand2_1 _21947_ (.A(_04344_),
    .B(_04345_),
    .Y(_04347_));
 sky130_fd_sc_hd__xnor2_1 _21948_ (.A(_04255_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_2 _21949_ (.A(net3670),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__o211ai_1 _21950_ (.A1(_04349_),
    .A2(_04250_),
    .B1(_08009_),
    .C1(net3756),
    .Y(_04350_));
 sky130_fd_sc_hd__nor2_1 _21951_ (.A(_10165_),
    .B(_10173_),
    .Y(_04351_));
 sky130_fd_sc_hd__xnor2_1 _21952_ (.A(net3726),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a221oi_1 _21953_ (.A1(_10165_),
    .A2(_10173_),
    .B1(_02127_),
    .B2(_04352_),
    .C1(_03273_),
    .Y(_04353_));
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(net3557),
    .B(_02391_),
    .Y(_04354_));
 sky130_fd_sc_hd__nor2_2 _21955_ (.A(_02182_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__mux2i_2 _21956_ (.A0(_03259_),
    .A1(_03262_),
    .S(net3619),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2b_1 _21957_ (.A_N(_04107_),
    .B(net3578),
    .Y(_04357_));
 sky130_fd_sc_hd__o211ai_1 _21958_ (.A1(net3578),
    .A2(_04356_),
    .B1(_04357_),
    .C1(net3558),
    .Y(_04358_));
 sky130_fd_sc_hd__o211ai_1 _21959_ (.A1(net3558),
    .A2(_02206_),
    .B1(_04358_),
    .C1(net3559),
    .Y(_04359_));
 sky130_fd_sc_hd__o211ai_1 _21960_ (.A1(net3559),
    .A2(_02705_),
    .B1(_04359_),
    .C1(net3560),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ai_4 _21961_ (.A1(net3560),
    .A2(_02404_),
    .B1(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _21962_ (.A(net3603),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__o21ai_0 _21963_ (.A1(_02057_),
    .A2(_04355_),
    .B1(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor4_1 _21964_ (.A(net3739),
    .B(net3738),
    .C(_04353_),
    .D(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__o21ai_4 _21965_ (.A1(net3486),
    .A2(_02702_),
    .B1(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__o21ai_4 _21966_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_13047_),
    .B1(_08501_),
    .Y(_04366_));
 sky130_fd_sc_hd__a21oi_4 _21967_ (.A1(_11473_),
    .A2(_04366_),
    .B1(net3472),
    .Y(_04367_));
 sky130_fd_sc_hd__mux4_2 _21968_ (.A0(net45),
    .A1(net28),
    .A2(net49),
    .A3(net36),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04368_));
 sky130_fd_sc_hd__nand2_1 _21969_ (.A(_01670_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__a21oi_2 _21970_ (.A1(_03086_),
    .A2(_04369_),
    .B1(net3469),
    .Y(_04370_));
 sky130_fd_sc_hd__a31oi_2 _21971_ (.A1(_04367_),
    .A2(_04365_),
    .A3(_04350_),
    .B1(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_405 ();
 sky130_fd_sc_hd__nand2_1 _21973_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .B(_02153_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21ai_0 _21974_ (.A1(_02153_),
    .A2(net3408),
    .B1(_04373_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2b_1 _21975_ (.A_N(_02529_),
    .B(net3670),
    .Y(_04374_));
 sky130_fd_sc_hd__nand2_1 _21976_ (.A(_04097_),
    .B(_04254_),
    .Y(_04375_));
 sky130_fd_sc_hd__inv_1 _21977_ (.A(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__and2_4 _21978_ (.A(_04251_),
    .B(_04344_),
    .X(_04377_));
 sky130_fd_sc_hd__a21bo_1 _21979_ (.A1(_04130_),
    .A2(_04376_),
    .B1_N(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__nor2_1 _21980_ (.A(_04258_),
    .B(_04341_),
    .Y(_04379_));
 sky130_fd_sc_hd__nand2_1 _21981_ (.A(_04258_),
    .B(_04341_),
    .Y(_04380_));
 sky130_fd_sc_hd__o21a_4 _21982_ (.A1(_04257_),
    .A2(_04379_),
    .B1(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__maj3_4 _21983_ (.A(_04303_),
    .B(_04320_),
    .C(_04340_),
    .X(_04382_));
 sky130_fd_sc_hd__o21ai_2 _21984_ (.A1(_04304_),
    .A2(_04317_),
    .B1(_04318_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21ai_0 _21985_ (.A1(_03460_),
    .A2(_04265_),
    .B1(_03459_),
    .Y(_04384_));
 sky130_fd_sc_hd__o21ai_2 _21986_ (.A1(net3627),
    .A2(_04269_),
    .B1(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__xor2_1 _21987_ (.A(_04299_),
    .B(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__xnor2_1 _21988_ (.A(_03803_),
    .B(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__maj3_4 _21989_ (.A(_03951_),
    .B(_04296_),
    .C(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _21990_ (.A(_02556_),
    .B(_03570_),
    .Y(_04389_));
 sky130_fd_sc_hd__nor2_1 _21991_ (.A(_02680_),
    .B(_02744_),
    .Y(_04390_));
 sky130_fd_sc_hd__nor2_2 _21992_ (.A(_02505_),
    .B(_02987_),
    .Y(_04391_));
 sky130_fd_sc_hd__xnor2_1 _21993_ (.A(_04390_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__xnor2_1 _21994_ (.A(_04389_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_2 _21995_ (.A(_02270_),
    .B(_02320_),
    .Y(_04394_));
 sky130_fd_sc_hd__a21oi_1 _21996_ (.A1(_04282_),
    .A2(_04394_),
    .B1(net3638),
    .Y(_04395_));
 sky130_fd_sc_hd__nor2_1 _21997_ (.A(_04282_),
    .B(_04286_),
    .Y(_04396_));
 sky130_fd_sc_hd__o21ai_2 _21998_ (.A1(_04395_),
    .A2(_04396_),
    .B1(net3630),
    .Y(_04397_));
 sky130_fd_sc_hd__xor2_1 _21999_ (.A(_04393_),
    .B(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__a21o_4 _22000_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net3668),
    .B1(net3732),
    .X(_04399_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_404 ();
 sky130_fd_sc_hd__a21oi_2 _22002_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_03681_),
    .B1(net3731),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _22003_ (.A(_03460_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__nor2_1 _22004_ (.A(_04269_),
    .B(_04299_),
    .Y(_04403_));
 sky130_fd_sc_hd__maj3_1 _22005_ (.A(net3629),
    .B(net3627),
    .C(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__nor2_1 _22006_ (.A(net3577),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__a21oi_1 _22007_ (.A1(_04269_),
    .A2(_04299_),
    .B1(_03460_),
    .Y(_04406_));
 sky130_fd_sc_hd__o22ai_1 _22008_ (.A1(_04265_),
    .A2(_04402_),
    .B1(_04406_),
    .B2(net3629),
    .Y(_04407_));
 sky130_fd_sc_hd__nor2_1 _22009_ (.A(_03803_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21o_4 _22010_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_03681_),
    .B1(net3731),
    .X(_04409_));
 sky130_fd_sc_hd__nand3_1 _22011_ (.A(net3629),
    .B(net3627),
    .C(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__o221ai_1 _22012_ (.A1(net3629),
    .A2(_04402_),
    .B1(_04405_),
    .B2(_04408_),
    .C1(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_2 _22013_ (.A(_04399_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__xor2_1 _22014_ (.A(_04290_),
    .B(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__xnor2_1 _22015_ (.A(_04398_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__xnor2_1 _22016_ (.A(_04388_),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__xnor2_1 _22017_ (.A(_04282_),
    .B(_04287_),
    .Y(_04416_));
 sky130_fd_sc_hd__maj3_1 _22018_ (.A(_04071_),
    .B(_04277_),
    .C(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nand2_2 _22019_ (.A(_04314_),
    .B(_04315_),
    .Y(_04418_));
 sky130_fd_sc_hd__or2_4 _22020_ (.A(net3633),
    .B(_02784_),
    .X(_04419_));
 sky130_fd_sc_hd__nand2b_2 _22021_ (.A_N(net3634),
    .B(_02859_),
    .Y(_04420_));
 sky130_fd_sc_hd__or3_4 _22022_ (.A(net471),
    .B(_08498_),
    .C(_10390_),
    .X(_04421_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_403 ();
 sky130_fd_sc_hd__nor2_4 _22024_ (.A(net3757),
    .B(_04421_),
    .Y(_04423_));
 sky130_fd_sc_hd__nand2_1 _22025_ (.A(_02476_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__xnor2_1 _22026_ (.A(_04420_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__xor2_1 _22027_ (.A(_04419_),
    .B(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__maj3_1 _22028_ (.A(_04306_),
    .B(_04307_),
    .C(_04308_),
    .X(_04427_));
 sky130_fd_sc_hd__maj3_1 _22029_ (.A(_04278_),
    .B(_04279_),
    .C(_04280_),
    .X(_04428_));
 sky130_fd_sc_hd__xnor2_1 _22030_ (.A(_04427_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__xnor2_1 _22031_ (.A(_04426_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__maj3_2 _22032_ (.A(_04311_),
    .B(_04310_),
    .C(_04312_),
    .X(_04431_));
 sky130_fd_sc_hd__xnor2_1 _22033_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__xor2_1 _22034_ (.A(_04418_),
    .B(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__xnor2_1 _22035_ (.A(_04417_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__xnor2_1 _22036_ (.A(_04415_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__xor2_1 _22037_ (.A(_04283_),
    .B(_04289_),
    .X(_04436_));
 sky130_fd_sc_hd__xnor2_1 _22038_ (.A(_03952_),
    .B(_04301_),
    .Y(_04437_));
 sky130_fd_sc_hd__maj3_1 _22039_ (.A(_04274_),
    .B(_04436_),
    .C(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__xnor2_1 _22040_ (.A(_04435_),
    .B(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__xor2_1 _22041_ (.A(_04383_),
    .B(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__xnor2_2 _22042_ (.A(_04382_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__nand2_2 _22043_ (.A(_04381_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__inv_1 _22044_ (.A(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__nor2_2 _22045_ (.A(_04381_),
    .B(_04441_),
    .Y(_04444_));
 sky130_fd_sc_hd__a211oi_1 _22046_ (.A1(_04345_),
    .A2(net3452),
    .B1(_04443_),
    .C1(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__o211a_1 _22047_ (.A1(_04443_),
    .A2(_04444_),
    .B1(_04345_),
    .C1(net3452),
    .X(_04446_));
 sky130_fd_sc_hd__o21ai_2 _22048_ (.A1(_04445_),
    .A2(_04446_),
    .B1(_02000_),
    .Y(_04447_));
 sky130_fd_sc_hd__a21oi_2 _22049_ (.A1(_04374_),
    .A2(_04447_),
    .B1(net3937),
    .Y(_04448_));
 sky130_fd_sc_hd__o21ai_0 _22050_ (.A1(_08009_),
    .A2(_10204_),
    .B1(net3756),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_1 _22051_ (.A(_10203_),
    .B(_10231_),
    .Y(_04450_));
 sky130_fd_sc_hd__xnor2_1 _22052_ (.A(_02133_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__o221ai_1 _22053_ (.A1(_10203_),
    .A2(_10231_),
    .B1(_02184_),
    .B2(_04451_),
    .C1(_02137_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand3_1 _22054_ (.A(net3746),
    .B(_11488_),
    .C(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__a221oi_2 _22055_ (.A1(net3602),
    .A2(_03254_),
    .B1(_03269_),
    .B2(net3603),
    .C1(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__o21ai_4 _22056_ (.A1(net3487),
    .A2(_02702_),
    .B1(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21a_4 _22057_ (.A1(_04448_),
    .A2(_04449_),
    .B1(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__mux4_2 _22058_ (.A0(net46),
    .A1(net29),
    .A2(net52),
    .A3(net37),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04457_));
 sky130_fd_sc_hd__nand2_1 _22059_ (.A(_01670_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand3_1 _22060_ (.A(net3472),
    .B(_03086_),
    .C(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__o21ai_2 _22061_ (.A1(net3472),
    .A2(_04456_),
    .B1(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_402 ();
 sky130_fd_sc_hd__nand2_1 _22063_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .B(_02153_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21ai_0 _22064_ (.A1(_02153_),
    .A2(net3407),
    .B1(_04462_),
    .Y(_00534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_401 ();
 sky130_fd_sc_hd__a22oi_1 _22066_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net48),
    .B1(_03238_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _22067_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_03772_),
    .Y(_04465_));
 sky130_fd_sc_hd__o21ai_0 _22068_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03771_),
    .B1(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__a221o_1 _22069_ (.A1(\load_store_unit_i.rdata_q[13] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[5] ),
    .C1(_02847_),
    .X(_04467_));
 sky130_fd_sc_hd__o21ai_2 _22070_ (.A1(_01670_),
    .A2(_04466_),
    .B1(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__o221ai_4 _22071_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03770_),
    .B1(_04464_),
    .B2(_03237_),
    .C1(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__nor2_4 _22072_ (.A(net3936),
    .B(_02225_),
    .Y(_04470_));
 sky130_fd_sc_hd__nor2_1 _22073_ (.A(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__a21oi_4 _22074_ (.A1(_03764_),
    .A2(_04470_),
    .B1(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__nand2_1 _22075_ (.A(net3625),
    .B(net3600),
    .Y(_04473_));
 sky130_fd_sc_hd__o21ai_0 _22076_ (.A1(_02184_),
    .A2(_04473_),
    .B1(_03272_),
    .Y(_04474_));
 sky130_fd_sc_hd__nand2_1 _22077_ (.A(_02133_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__o21ai_0 _22078_ (.A1(net3625),
    .A2(net3600),
    .B1(_02133_),
    .Y(_04476_));
 sky130_fd_sc_hd__nand2_1 _22079_ (.A(_04473_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__a22oi_1 _22080_ (.A1(net3602),
    .A2(_04361_),
    .B1(_04475_),
    .B2(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21ai_2 _22081_ (.A1(_02020_),
    .A2(_04355_),
    .B1(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__a211o_4 _22082_ (.A1(net3537),
    .A2(_02006_),
    .B1(_04479_),
    .C1(net3755),
    .X(_04480_));
 sky130_fd_sc_hd__o21ai_4 _22083_ (.A1(net3747),
    .A2(_04472_),
    .B1(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand3_4 _22084_ (.A(_11645_),
    .B(_01655_),
    .C(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__o21ai_4 _22085_ (.A1(net3469),
    .A2(_04469_),
    .B1(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_400 ();
 sky130_fd_sc_hd__nand2_1 _22087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .B(_03280_),
    .Y(_04485_));
 sky130_fd_sc_hd__o21ai_0 _22088_ (.A1(_03280_),
    .A2(_04483_),
    .B1(_04485_),
    .Y(_00535_));
 sky130_fd_sc_hd__inv_1 _22089_ (.A(_04345_),
    .Y(_04486_));
 sky130_fd_sc_hd__a21boi_0 _22090_ (.A1(_04252_),
    .A2(_04376_),
    .B1_N(_04377_),
    .Y(_04487_));
 sky130_fd_sc_hd__o31ai_1 _22091_ (.A1(_04486_),
    .A2(_04444_),
    .A3(_04487_),
    .B1(_04442_),
    .Y(_04488_));
 sky130_fd_sc_hd__inv_1 _22092_ (.A(_04439_),
    .Y(_04489_));
 sky130_fd_sc_hd__maj3_4 _22093_ (.A(_04382_),
    .B(_04383_),
    .C(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_399 ();
 sky130_fd_sc_hd__xnor2_1 _22095_ (.A(net3571),
    .B(_04412_),
    .Y(_04492_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_397 ();
 sky130_fd_sc_hd__o22ai_1 _22098_ (.A1(_03460_),
    .A2(_04299_),
    .B1(_04402_),
    .B2(_04169_),
    .Y(_04495_));
 sky130_fd_sc_hd__nand2_1 _22099_ (.A(net3629),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_395 ();
 sky130_fd_sc_hd__nand4_1 _22102_ (.A(_03459_),
    .B(net3627),
    .C(_04265_),
    .D(_04401_),
    .Y(_04499_));
 sky130_fd_sc_hd__a21oi_1 _22103_ (.A1(_04496_),
    .A2(_04499_),
    .B1(_04399_),
    .Y(_04500_));
 sky130_fd_sc_hd__a21oi_2 _22104_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(_03681_),
    .B1(net3731),
    .Y(_04501_));
 sky130_fd_sc_hd__o21ai_0 _22105_ (.A1(_03460_),
    .A2(_04409_),
    .B1(_03459_),
    .Y(_04502_));
 sky130_fd_sc_hd__o21ai_0 _22106_ (.A1(net3627),
    .A2(_04299_),
    .B1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand3_1 _22107_ (.A(_04409_),
    .B(_04385_),
    .C(_04501_),
    .Y(_04504_));
 sky130_fd_sc_hd__o211ai_1 _22108_ (.A1(_04501_),
    .A2(_04503_),
    .B1(_04504_),
    .C1(_03803_),
    .Y(_04505_));
 sky130_fd_sc_hd__o21ai_2 _22109_ (.A1(_03803_),
    .A2(_04500_),
    .B1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__o21ai_2 _22110_ (.A1(_03951_),
    .A2(_04492_),
    .B1(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__nand2_2 _22111_ (.A(_02900_),
    .B(_03570_),
    .Y(_04508_));
 sky130_fd_sc_hd__xnor2_1 _22112_ (.A(_02505_),
    .B(_02556_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _22113_ (.A(net3630),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__xnor2_1 _22114_ (.A(_04508_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__a21oi_1 _22115_ (.A1(_04393_),
    .A2(_04394_),
    .B1(net3638),
    .Y(_04512_));
 sky130_fd_sc_hd__nor2_1 _22116_ (.A(_04286_),
    .B(_04393_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_1 _22117_ (.A1(_04512_),
    .A2(_04513_),
    .B1(net3630),
    .Y(_04514_));
 sky130_fd_sc_hd__xor2_1 _22118_ (.A(_04511_),
    .B(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_394 ();
 sky130_fd_sc_hd__a21oi_4 _22120_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net3668),
    .B1(net3732),
    .Y(_04517_));
 sky130_fd_sc_hd__nor2_1 _22121_ (.A(net3628),
    .B(_04399_),
    .Y(_04518_));
 sky130_fd_sc_hd__o21ai_0 _22122_ (.A1(_04409_),
    .A2(_04399_),
    .B1(net3628),
    .Y(_04519_));
 sky130_fd_sc_hd__a22oi_1 _22123_ (.A1(_04401_),
    .A2(_04518_),
    .B1(_04519_),
    .B2(_03459_),
    .Y(_04520_));
 sky130_fd_sc_hd__nor2_1 _22124_ (.A(_03460_),
    .B(_04501_),
    .Y(_04521_));
 sky130_fd_sc_hd__o21ai_0 _22125_ (.A1(_04401_),
    .A2(_04501_),
    .B1(_03460_),
    .Y(_04522_));
 sky130_fd_sc_hd__a221oi_1 _22126_ (.A1(_04409_),
    .A2(_04521_),
    .B1(_04522_),
    .B2(net3629),
    .C1(_03691_),
    .Y(_04523_));
 sky130_fd_sc_hd__a21oi_1 _22127_ (.A1(net3577),
    .A2(_04520_),
    .B1(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand2_1 _22128_ (.A(net3628),
    .B(_04399_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _22129_ (.A(_03459_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a211oi_1 _22130_ (.A1(_03459_),
    .A2(_04518_),
    .B1(_04524_),
    .C1(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__xnor2_2 _22131_ (.A(_04517_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__xnor2_1 _22132_ (.A(_04290_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__xnor2_1 _22133_ (.A(_04515_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__xnor2_1 _22134_ (.A(_04507_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2_2 _22135_ (.A(_04430_),
    .B(_04431_),
    .Y(_04532_));
 sky130_fd_sc_hd__maj3_1 _22136_ (.A(_04419_),
    .B(_04420_),
    .C(_04424_),
    .X(_04533_));
 sky130_fd_sc_hd__nor2_1 _22137_ (.A(_02744_),
    .B(net3632),
    .Y(_04534_));
 sky130_fd_sc_hd__nor2_1 _22138_ (.A(net3633),
    .B(_02856_),
    .Y(_04535_));
 sky130_fd_sc_hd__and3_4 _22139_ (.A(net3760),
    .B(net3634),
    .C(_03058_),
    .X(_04536_));
 sky130_fd_sc_hd__xor2_1 _22140_ (.A(_04535_),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__xnor2_1 _22141_ (.A(_04534_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__o22ai_1 _22142_ (.A1(_02680_),
    .A2(_02744_),
    .B1(_02877_),
    .B2(_02764_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor4_1 _22143_ (.A(_02764_),
    .B(_02680_),
    .C(_02744_),
    .D(_02877_),
    .Y(_04540_));
 sky130_fd_sc_hd__a21oi_2 _22144_ (.A1(_04391_),
    .A2(_04539_),
    .B1(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__xnor2_1 _22145_ (.A(_04538_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__xnor2_1 _22146_ (.A(_04533_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__maj3_1 _22147_ (.A(_04427_),
    .B(_04426_),
    .C(_04428_),
    .X(_04544_));
 sky130_fd_sc_hd__xor2_1 _22148_ (.A(_04543_),
    .B(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__xor2_1 _22149_ (.A(_04532_),
    .B(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__xnor2_1 _22150_ (.A(_04287_),
    .B(_04393_),
    .Y(_04547_));
 sky130_fd_sc_hd__maj3_4 _22151_ (.A(_04071_),
    .B(_04397_),
    .C(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__xnor2_2 _22152_ (.A(_04546_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__xnor2_1 _22153_ (.A(_04531_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__xnor2_1 _22154_ (.A(_04289_),
    .B(_04398_),
    .Y(_04551_));
 sky130_fd_sc_hd__xnor2_1 _22155_ (.A(_03952_),
    .B(_04412_),
    .Y(_04552_));
 sky130_fd_sc_hd__maj3_1 _22156_ (.A(_04388_),
    .B(_04551_),
    .C(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _22157_ (.A(_04550_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__maj3_4 _22158_ (.A(_04418_),
    .B(_04417_),
    .C(_04432_),
    .X(_04555_));
 sky130_fd_sc_hd__nor2_1 _22159_ (.A(_04415_),
    .B(_04434_),
    .Y(_04556_));
 sky130_fd_sc_hd__nand2_1 _22160_ (.A(_04415_),
    .B(_04434_),
    .Y(_04557_));
 sky130_fd_sc_hd__o21ai_2 _22161_ (.A1(_04556_),
    .A2(_04438_),
    .B1(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__xnor2_1 _22162_ (.A(_04555_),
    .B(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__xnor2_2 _22163_ (.A(_04554_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nor2_2 _22164_ (.A(_04490_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2_2 _22165_ (.A(_04490_),
    .B(_04560_),
    .Y(_04562_));
 sky130_fd_sc_hd__nor2b_1 _22166_ (.A(_04561_),
    .B_N(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__xor2_1 _22167_ (.A(_04563_),
    .B(_04488_),
    .X(_04564_));
 sky130_fd_sc_hd__mux2i_2 _22168_ (.A0(_02605_),
    .A1(_04564_),
    .S(_02000_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _22169_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .Y(_04566_));
 sky130_fd_sc_hd__o21ai_4 _22170_ (.A1(_04565_),
    .A2(net3937),
    .B1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__mux4_2 _22171_ (.A0(net47),
    .A1(net30),
    .A2(net53),
    .A3(net39),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04568_));
 sky130_fd_sc_hd__a21oi_4 _22172_ (.A1(_01670_),
    .A2(_04568_),
    .B1(_03289_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _22173_ (.A(net321),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor2_1 _22174_ (.A(_10269_),
    .B(_02020_),
    .Y(_04571_));
 sky130_fd_sc_hd__nor2_1 _22175_ (.A(net3599),
    .B(net3603),
    .Y(_04572_));
 sky130_fd_sc_hd__nor2_1 _22176_ (.A(_04571_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__mux2i_1 _22177_ (.A0(_03257_),
    .A1(_04573_),
    .S(net3621),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2b_1 _22178_ (.A_N(_04356_),
    .B(net3578),
    .Y(_04575_));
 sky130_fd_sc_hd__o211ai_1 _22179_ (.A1(net3578),
    .A2(_04574_),
    .B1(_04575_),
    .C1(net3558),
    .Y(_04576_));
 sky130_fd_sc_hd__o21ai_0 _22180_ (.A1(net3558),
    .A2(_04108_),
    .B1(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__nand2_1 _22181_ (.A(net3559),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__o21ai_1 _22182_ (.A1(net3559),
    .A2(_02450_),
    .B1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor2_1 _22183_ (.A(net3560),
    .B(_02616_),
    .Y(_04580_));
 sky130_fd_sc_hd__a21o_4 _22184_ (.A1(net3560),
    .A2(_04579_),
    .B1(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _22185_ (.A(net3603),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_2 _22186_ (.A(_02171_),
    .B(_02056_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _22187_ (.A(_02435_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_4 _22188_ (.A1(_02077_),
    .A2(_04583_),
    .B1(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nor2_1 _22189_ (.A(_10269_),
    .B(_10296_),
    .Y(_04586_));
 sky130_fd_sc_hd__xnor2_1 _22190_ (.A(_02133_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a221oi_1 _22191_ (.A1(_10269_),
    .A2(_10296_),
    .B1(_02127_),
    .B2(_04587_),
    .C1(_03273_),
    .Y(_04588_));
 sky130_fd_sc_hd__a21oi_1 _22192_ (.A1(net3602),
    .A2(_04585_),
    .B1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__o211ai_1 _22193_ (.A1(net3485),
    .A2(_02702_),
    .B1(_04582_),
    .C1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_2 _22194_ (.A(net3744),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a31oi_4 _22195_ (.A1(_11503_),
    .A2(_01655_),
    .A3(_04591_),
    .B1(_04569_),
    .Y(_04592_));
 sky130_fd_sc_hd__a21oi_2 _22196_ (.A1(_04567_),
    .A2(_04570_),
    .B1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_393 ();
 sky130_fd_sc_hd__nand2_1 _22198_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .B(_02153_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_0 _22199_ (.A1(_02153_),
    .A2(net3406),
    .B1(_04595_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _22200_ (.A(_04345_),
    .B(_04378_),
    .Y(_04596_));
 sky130_fd_sc_hd__and2_4 _22201_ (.A(_04442_),
    .B(_04562_),
    .X(_04597_));
 sky130_fd_sc_hd__and2_4 _22202_ (.A(_04444_),
    .B(_04562_),
    .X(_04598_));
 sky130_fd_sc_hd__a211oi_2 _22203_ (.A1(_04596_),
    .A2(_04597_),
    .B1(_04598_),
    .C1(_04561_),
    .Y(_04599_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_04555_),
    .B(_04554_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2_1 _22205_ (.A(_04555_),
    .B(_04554_),
    .Y(_04601_));
 sky130_fd_sc_hd__o21ai_2 _22206_ (.A1(_04558_),
    .A2(_04600_),
    .B1(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _22207_ (.A(_04531_),
    .B(_04549_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2_1 _22208_ (.A(_04603_),
    .B(_04553_),
    .Y(_04604_));
 sky130_fd_sc_hd__o21ai_2 _22209_ (.A1(_04531_),
    .A2(_04549_),
    .B1(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__xor2_1 _22210_ (.A(_04289_),
    .B(_04515_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_2 _22211_ (.A(net3571),
    .B(net3570),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_4 _22212_ (.A(_04039_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__xnor2_1 _22213_ (.A(_04608_),
    .B(_04528_),
    .Y(_04609_));
 sky130_fd_sc_hd__maj3_1 _22214_ (.A(_04507_),
    .B(_04606_),
    .C(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__nor2b_4 _22215_ (.A(_04543_),
    .B_N(_04544_),
    .Y(_04611_));
 sky130_fd_sc_hd__xnor2_1 _22216_ (.A(_04287_),
    .B(_04511_),
    .Y(_04612_));
 sky130_fd_sc_hd__maj3_2 _22217_ (.A(_04071_),
    .B(_04514_),
    .C(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__nor2_2 _22218_ (.A(net3632),
    .B(_02877_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_2 _22219_ (.A(_02744_),
    .B(_02856_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_1 _22220_ (.A(net3633),
    .B(_04423_),
    .Y(_04616_));
 sky130_fd_sc_hd__xnor2_1 _22221_ (.A(_04615_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__xnor2_1 _22222_ (.A(_04614_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__maj3_1 _22223_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .X(_04619_));
 sky130_fd_sc_hd__maj3_1 _22224_ (.A(_02505_),
    .B(_02764_),
    .C(_04508_),
    .X(_04620_));
 sky130_fd_sc_hd__nand2b_4 _22225_ (.A_N(_04620_),
    .B(net3630),
    .Y(_04621_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_392 ();
 sky130_fd_sc_hd__xnor2_1 _22227_ (.A(_04619_),
    .B(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__xnor2_1 _22228_ (.A(_04618_),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__maj3_1 _22229_ (.A(_04533_),
    .B(_04538_),
    .C(_04541_),
    .X(_04625_));
 sky130_fd_sc_hd__inv_1 _22230_ (.A(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__xnor2_1 _22231_ (.A(_04624_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__xnor3_1 _22232_ (.A(_04611_),
    .B(_04613_),
    .C(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_391 ();
 sky130_fd_sc_hd__nor3_1 _22234_ (.A(net3627),
    .B(_04401_),
    .C(_04399_),
    .Y(_04630_));
 sky130_fd_sc_hd__o21ai_0 _22235_ (.A1(_04521_),
    .A2(_04630_),
    .B1(net3629),
    .Y(_04631_));
 sky130_fd_sc_hd__o31ai_1 _22236_ (.A1(_03470_),
    .A2(_04401_),
    .A3(_04399_),
    .B1(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ai_0 _22237_ (.A1(_03460_),
    .A2(_04399_),
    .B1(_03459_),
    .Y(_04633_));
 sky130_fd_sc_hd__o21ai_2 _22238_ (.A1(net3628),
    .A2(_04501_),
    .B1(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor2_1 _22239_ (.A(_04517_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__a31oi_1 _22240_ (.A1(_04399_),
    .A2(_04503_),
    .A3(_04517_),
    .B1(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__nor2_1 _22241_ (.A(net3577),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__a31oi_2 _22242_ (.A1(net3577),
    .A2(_04517_),
    .A3(_04632_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__xnor2_1 _22243_ (.A(_03951_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__a21o_1 _22244_ (.A1(_04038_),
    .A2(_03951_),
    .B1(_04638_),
    .X(_04640_));
 sky130_fd_sc_hd__o21ai_0 _22245_ (.A1(_03951_),
    .A2(_04528_),
    .B1(_04638_),
    .Y(_04641_));
 sky130_fd_sc_hd__a22oi_1 _22246_ (.A1(net3571),
    .A2(_04639_),
    .B1(_04640_),
    .B2(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2_1 _22247_ (.A(_02680_),
    .B(_04287_),
    .Y(_04643_));
 sky130_fd_sc_hd__o21ai_1 _22248_ (.A1(_04287_),
    .A2(_04508_),
    .B1(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__xnor2_2 _22249_ (.A(_04509_),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_8 _22250_ (.A(net3630),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__a21oi_1 _22251_ (.A1(_04394_),
    .A2(_04511_),
    .B1(net3638),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_1 _22252_ (.A(_04286_),
    .B(_04511_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_2 _22253_ (.A1(_04647_),
    .A2(_04648_),
    .B1(net3630),
    .Y(_04649_));
 sky130_fd_sc_hd__xnor2_2 _22254_ (.A(_04072_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__xnor2_4 _22255_ (.A(_04646_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__a21o_4 _22256_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net3668),
    .B1(net3732),
    .X(_04652_));
 sky130_fd_sc_hd__nor2_1 _22257_ (.A(_03460_),
    .B(_04517_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _22258_ (.A(net3629),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_390 ();
 sky130_fd_sc_hd__nand3_1 _22260_ (.A(_03459_),
    .B(_03460_),
    .C(_04517_),
    .Y(_04656_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_389 ();
 sky130_fd_sc_hd__a21o_4 _22262_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net3668),
    .B1(net3732),
    .X(_04658_));
 sky130_fd_sc_hd__a21oi_1 _22263_ (.A1(_04399_),
    .A2(_04658_),
    .B1(net3628),
    .Y(_04659_));
 sky130_fd_sc_hd__o22ai_1 _22264_ (.A1(_04517_),
    .A2(_04525_),
    .B1(_04659_),
    .B2(_03459_),
    .Y(_04660_));
 sky130_fd_sc_hd__o21ai_0 _22265_ (.A1(_04399_),
    .A2(_04658_),
    .B1(net3628),
    .Y(_04661_));
 sky130_fd_sc_hd__a221o_1 _22266_ (.A1(_04517_),
    .A2(_04518_),
    .B1(_04661_),
    .B2(_03459_),
    .C1(_03803_),
    .X(_04662_));
 sky130_fd_sc_hd__o21ai_1 _22267_ (.A1(net3577),
    .A2(_04660_),
    .B1(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand3_2 _22268_ (.A(_04654_),
    .B(_04656_),
    .C(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__xnor2_4 _22269_ (.A(_04652_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__xnor2_1 _22270_ (.A(_04651_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__xnor2_1 _22271_ (.A(_04642_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__xor2_1 _22272_ (.A(_04628_),
    .B(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__xnor2_1 _22273_ (.A(_04610_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__maj3_4 _22274_ (.A(_04532_),
    .B(_04545_),
    .C(_04548_),
    .X(_04670_));
 sky130_fd_sc_hd__xnor2_1 _22275_ (.A(_04669_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_1 _22276_ (.A(_04605_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__or2_4 _22277_ (.A(_04602_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__nand2_2 _22278_ (.A(_04602_),
    .B(_04672_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _22279_ (.A(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xor2_1 _22280_ (.A(_04599_),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_2 _22281_ (.A(_02000_),
    .B(_02698_),
    .Y(_04677_));
 sky130_fd_sc_hd__a211oi_4 _22282_ (.A1(_02000_),
    .A2(_04676_),
    .B1(_04677_),
    .C1(net3937),
    .Y(_04678_));
 sky130_fd_sc_hd__and2_0 _22283_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _22284_ (.A(net3474),
    .B(_02006_),
    .Y(_04680_));
 sky130_fd_sc_hd__nor2_1 _22285_ (.A(_10336_),
    .B(_02020_),
    .Y(_04681_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(net3598),
    .B(net3603),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _22287_ (.A(_04681_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__nor2_1 _22288_ (.A(net3619),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(net3621),
    .B(_04573_),
    .Y(_04685_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(_04684_),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _22291_ (.A(net3578),
    .B(_03260_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21ai_0 _22292_ (.A1(net3578),
    .A2(_04686_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_1 _22293_ (.A(net3558),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__o211ai_1 _22294_ (.A1(net3558),
    .A2(_04226_),
    .B1(_04689_),
    .C1(_02016_),
    .Y(_04690_));
 sky130_fd_sc_hd__o211ai_1 _22295_ (.A1(_02016_),
    .A2(_02395_),
    .B1(_04690_),
    .C1(net3560),
    .Y(_04691_));
 sky130_fd_sc_hd__o21ai_4 _22296_ (.A1(net3560),
    .A2(_02714_),
    .B1(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21ai_4 _22297_ (.A1(_02171_),
    .A2(_02710_),
    .B1(_02612_),
    .Y(_04693_));
 sky130_fd_sc_hd__nor2_1 _22298_ (.A(_10336_),
    .B(_10366_),
    .Y(_04694_));
 sky130_fd_sc_hd__xor2_1 _22299_ (.A(_02133_),
    .B(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__nand2_1 _22300_ (.A(_10336_),
    .B(_10366_),
    .Y(_04696_));
 sky130_fd_sc_hd__o211ai_1 _22301_ (.A1(_02184_),
    .A2(_04695_),
    .B1(_04696_),
    .C1(_02137_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand3_1 _22302_ (.A(net3746),
    .B(_11527_),
    .C(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__a221oi_4 _22303_ (.A1(net3603),
    .A2(_04692_),
    .B1(_04693_),
    .B2(net3602),
    .C1(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_4 _22304_ (.A1(_04680_),
    .A2(_04699_),
    .B1(net3472),
    .Y(_04700_));
 sky130_fd_sc_hd__o21ai_2 _22305_ (.A1(_04678_),
    .A2(_04679_),
    .B1(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_388 ();
 sky130_fd_sc_hd__mux4_2 _22307_ (.A0(net48),
    .A1(net31),
    .A2(net54),
    .A3(net40),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04703_));
 sky130_fd_sc_hd__nand2_1 _22308_ (.A(_01670_),
    .B(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_1 _22309_ (.A1(_03086_),
    .A2(_04704_),
    .B1(net3469),
    .Y(_04705_));
 sky130_fd_sc_hd__a21oi_2 _22310_ (.A1(net3743),
    .A2(_04700_),
    .B1(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_387 ();
 sky130_fd_sc_hd__nor2_1 _22312_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .B(_03095_),
    .Y(_04708_));
 sky130_fd_sc_hd__a31oi_1 _22313_ (.A1(_03095_),
    .A2(net3405),
    .A3(net3457),
    .B1(_04708_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _22314_ (.A(net480),
    .B(_02006_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(_10452_),
    .B(_02020_),
    .Y(_04710_));
 sky130_fd_sc_hd__a21oi_1 _22316_ (.A1(net3597),
    .A2(_02020_),
    .B1(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__mux2i_1 _22317_ (.A0(_04683_),
    .A1(_04711_),
    .S(net3621),
    .Y(_04712_));
 sky130_fd_sc_hd__mux4_2 _22318_ (.A0(_04356_),
    .A1(_04712_),
    .A2(_04107_),
    .A3(_04574_),
    .S0(_02051_),
    .S1(net3578),
    .X(_04713_));
 sky130_fd_sc_hd__nand2_1 _22319_ (.A(_02056_),
    .B(_02208_),
    .Y(_04714_));
 sky130_fd_sc_hd__o211ai_1 _22320_ (.A1(_02056_),
    .A2(_04713_),
    .B1(_04714_),
    .C1(net3560),
    .Y(_04715_));
 sky130_fd_sc_hd__o21ai_4 _22321_ (.A1(net3560),
    .A2(_02820_),
    .B1(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__o21ai_2 _22322_ (.A1(_02171_),
    .A2(_02822_),
    .B1(_02612_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _22323_ (.A(net3602),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21ai_2 _22324_ (.A1(net3666),
    .A2(_10450_),
    .B1(_10451_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _22325_ (.A(_04719_),
    .B(_10480_),
    .Y(_04720_));
 sky130_fd_sc_hd__xnor2_1 _22326_ (.A(_02133_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o221ai_1 _22327_ (.A1(_04719_),
    .A2(_10480_),
    .B1(_02184_),
    .B2(_04721_),
    .C1(_02137_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _22328_ (.A(_04718_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__a21oi_4 _22329_ (.A1(net3603),
    .A2(_04716_),
    .B1(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__o21ai_2 _22330_ (.A1(_04490_),
    .A2(_04560_),
    .B1(_04674_),
    .Y(_04725_));
 sky130_fd_sc_hd__o21ai_0 _22331_ (.A1(_04486_),
    .A2(_04444_),
    .B1(_04597_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2b_1 _22332_ (.A_N(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__or3_1 _22333_ (.A(_03780_),
    .B(_04007_),
    .C(_04375_),
    .X(_04728_));
 sky130_fd_sc_hd__a21o_1 _22334_ (.A1(_04013_),
    .A2(_04099_),
    .B1(_04375_),
    .X(_04729_));
 sky130_fd_sc_hd__o2111a_1 _22335_ (.A1(_03779_),
    .A2(_04728_),
    .B1(_04729_),
    .C1(_04377_),
    .D1(_04597_),
    .X(_04730_));
 sky130_fd_sc_hd__o21ai_1 _22336_ (.A1(_04727_),
    .A2(_04730_),
    .B1(_04673_),
    .Y(_04731_));
 sky130_fd_sc_hd__maj3_4 _22337_ (.A(_04605_),
    .B(_04669_),
    .C(_04670_),
    .X(_04732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_386 ();
 sky130_fd_sc_hd__xnor2_1 _22339_ (.A(_04608_),
    .B(_04665_),
    .Y(_04734_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_384 ();
 sky130_fd_sc_hd__nand3b_1 _22342_ (.A_N(_04665_),
    .B(_04528_),
    .C(net3571),
    .Y(_04737_));
 sky130_fd_sc_hd__or3b_1 _22343_ (.A(net3571),
    .B(_04528_),
    .C_N(_04665_),
    .X(_04738_));
 sky130_fd_sc_hd__xor2_4 _22344_ (.A(_04646_),
    .B(_04650_),
    .X(_04739_));
 sky130_fd_sc_hd__nor2_1 _22345_ (.A(net3570),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__a31oi_1 _22346_ (.A1(net3570),
    .A2(_04737_),
    .A3(_04738_),
    .B1(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__o22a_1 _22347_ (.A1(_04528_),
    .A2(_04651_),
    .B1(_04665_),
    .B2(net3570),
    .X(_04742_));
 sky130_fd_sc_hd__a221oi_1 _22348_ (.A1(_04528_),
    .A2(_04739_),
    .B1(_04665_),
    .B2(_03951_),
    .C1(_04038_),
    .Y(_04743_));
 sky130_fd_sc_hd__a21oi_1 _22349_ (.A1(_04038_),
    .A2(_04742_),
    .B1(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__o21ai_0 _22350_ (.A1(_04741_),
    .A2(_04744_),
    .B1(_04638_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21ai_2 _22351_ (.A1(_04651_),
    .A2(_04734_),
    .B1(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__maj3_4 _22352_ (.A(_04071_),
    .B(_04646_),
    .C(_04649_),
    .X(_04747_));
 sky130_fd_sc_hd__nand2_1 _22353_ (.A(_04624_),
    .B(_04626_),
    .Y(_04748_));
 sky130_fd_sc_hd__inv_1 _22354_ (.A(_04619_),
    .Y(_04749_));
 sky130_fd_sc_hd__maj3_1 _22355_ (.A(_04618_),
    .B(_04749_),
    .C(_04621_),
    .X(_04750_));
 sky130_fd_sc_hd__nor2_2 _22356_ (.A(net3632),
    .B(_02987_),
    .Y(_04751_));
 sky130_fd_sc_hd__nor2_2 _22357_ (.A(_02856_),
    .B(_02877_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_2 _22358_ (.A(_02744_),
    .B(_03181_),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_1 _22359_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__xnor2_1 _22360_ (.A(_04751_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_04614_),
    .B(_04615_),
    .Y(_04756_));
 sky130_fd_sc_hd__nor2_1 _22362_ (.A(_04616_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__a21oi_2 _22363_ (.A1(_04614_),
    .A2(_04615_),
    .B1(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__xnor2_1 _22364_ (.A(_04621_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__xnor2_1 _22365_ (.A(_04755_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__xnor2_1 _22366_ (.A(_04750_),
    .B(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__xor2_1 _22367_ (.A(_04748_),
    .B(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__xnor2_1 _22368_ (.A(_04747_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_383 ();
 sky130_fd_sc_hd__a21oi_4 _22370_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net3668),
    .B1(net3732),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _22371_ (.A(_04399_),
    .B(_04517_),
    .Y(_04766_));
 sky130_fd_sc_hd__nor2_1 _22372_ (.A(net3628),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__o21ai_0 _22373_ (.A1(_04653_),
    .A2(_04767_),
    .B1(net3629),
    .Y(_04768_));
 sky130_fd_sc_hd__o21ai_2 _22374_ (.A1(_03470_),
    .A2(_04766_),
    .B1(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21ai_0 _22375_ (.A1(net3627),
    .A2(_04517_),
    .B1(net3629),
    .Y(_04770_));
 sky130_fd_sc_hd__o21ai_0 _22376_ (.A1(_03460_),
    .A2(_04658_),
    .B1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_1 _22377_ (.A(_04652_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand3_1 _22378_ (.A(_04658_),
    .B(_04634_),
    .C(_04765_),
    .Y(_04773_));
 sky130_fd_sc_hd__a21oi_2 _22379_ (.A1(_04772_),
    .A2(_04773_),
    .B1(net3577),
    .Y(_04774_));
 sky130_fd_sc_hd__a31oi_4 _22380_ (.A1(net3577),
    .A2(_04765_),
    .A3(_04769_),
    .B1(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__nor2_1 _22381_ (.A(net3570),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__xnor2_1 _22382_ (.A(net3570),
    .B(_04775_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand3_1 _22383_ (.A(net3570),
    .B(_04665_),
    .C(_04775_),
    .Y(_04778_));
 sky130_fd_sc_hd__o21ai_0 _22384_ (.A1(net3571),
    .A2(_04777_),
    .B1(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__a21oi_1 _22385_ (.A1(net3571),
    .A2(_04776_),
    .B1(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21oi_4 _22386_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(_10746_),
    .B1(net3669),
    .Y(_04781_));
 sky130_fd_sc_hd__nor3_1 _22387_ (.A(_03459_),
    .B(_03460_),
    .C(_04765_),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_1 _22388_ (.A(_03460_),
    .B(_04765_),
    .Y(_04783_));
 sky130_fd_sc_hd__o21ai_0 _22389_ (.A1(_04517_),
    .A2(_04765_),
    .B1(_03460_),
    .Y(_04784_));
 sky130_fd_sc_hd__a22oi_1 _22390_ (.A1(_04658_),
    .A2(_04783_),
    .B1(_04784_),
    .B2(net3629),
    .Y(_04785_));
 sky130_fd_sc_hd__nor2_1 _22391_ (.A(net3577),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__nor2_1 _22392_ (.A(net3628),
    .B(_04652_),
    .Y(_04787_));
 sky130_fd_sc_hd__o21ai_0 _22393_ (.A1(_04658_),
    .A2(_04652_),
    .B1(net3628),
    .Y(_04788_));
 sky130_fd_sc_hd__a22oi_1 _22394_ (.A1(_04517_),
    .A2(_04787_),
    .B1(_04788_),
    .B2(_03459_),
    .Y(_04789_));
 sky130_fd_sc_hd__nor2_1 _22395_ (.A(_03803_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__a2111oi_0 _22396_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(_10746_),
    .B1(net3629),
    .C1(net3627),
    .D1(net3669),
    .Y(_04791_));
 sky130_fd_sc_hd__nor4_1 _22397_ (.A(_04782_),
    .B(_04786_),
    .C(_04790_),
    .D(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__xnor2_1 _22398_ (.A(_04781_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__xnor2_1 _22399_ (.A(_04651_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__xnor2_1 _22400_ (.A(_04780_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__xnor2_1 _22401_ (.A(_04763_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__xor2_1 _22402_ (.A(_04746_),
    .B(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__nand2_1 _22403_ (.A(_04613_),
    .B(_04627_),
    .Y(_04798_));
 sky130_fd_sc_hd__nor2_1 _22404_ (.A(_04613_),
    .B(_04627_),
    .Y(_04799_));
 sky130_fd_sc_hd__a21oi_2 _22405_ (.A1(_04611_),
    .A2(_04798_),
    .B1(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _22406_ (.A(_04628_),
    .B(_04667_),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _22407_ (.A(_04628_),
    .B(_04667_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_1 _22408_ (.A1(_04610_),
    .A2(_04801_),
    .B1(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__nor2_2 _22409_ (.A(_04800_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2_1 _22410_ (.A(_04800_),
    .B(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2b_2 _22411_ (.A(_04804_),
    .B_N(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__xnor2_2 _22412_ (.A(_04797_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__nor2_2 _22413_ (.A(_04732_),
    .B(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand2_2 _22414_ (.A(_04732_),
    .B(_04807_),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2b_1 _22415_ (.A(_04808_),
    .B_N(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__xnor2_1 _22416_ (.A(_04731_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__mux2i_4 _22417_ (.A0(_02814_),
    .A1(_04811_),
    .S(_02000_),
    .Y(_04812_));
 sky130_fd_sc_hd__mux2i_4 _22418_ (.A0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A1(_04812_),
    .S(_08009_),
    .Y(_04813_));
 sky130_fd_sc_hd__a32o_1 _22419_ (.A1(_08498_),
    .A2(_04709_),
    .A3(_04724_),
    .B1(_04813_),
    .B2(net3756),
    .X(_04814_));
 sky130_fd_sc_hd__mux4_2 _22420_ (.A0(net50),
    .A1(net32),
    .A2(net55),
    .A3(net41),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04815_));
 sky130_fd_sc_hd__a21oi_2 _22421_ (.A1(_01670_),
    .A2(_04815_),
    .B1(_03289_),
    .Y(_04816_));
 sky130_fd_sc_hd__a31oi_2 _22422_ (.A1(_11548_),
    .A2(net3469),
    .A3(_04814_),
    .B1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_382 ();
 sky130_fd_sc_hd__mux2_1 _22424_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .A1(net3404),
    .S(_03095_),
    .X(_00538_));
 sky130_fd_sc_hd__maj3_2 _22425_ (.A(_04748_),
    .B(_04747_),
    .C(_04761_),
    .X(_04819_));
 sky130_fd_sc_hd__a21oi_4 _22426_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net3668),
    .B1(net3732),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _22427_ (.A(_03803_),
    .B(_04785_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _22428_ (.A(net3577),
    .B(_04789_),
    .Y(_04822_));
 sky130_fd_sc_hd__a221o_1 _22429_ (.A1(_03459_),
    .A2(_04787_),
    .B1(_04821_),
    .B2(_04822_),
    .C1(_04782_),
    .X(_04823_));
 sky130_fd_sc_hd__xnor2_2 _22430_ (.A(_04820_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__and3_1 _22431_ (.A(net3571),
    .B(_04665_),
    .C(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__nor3_1 _22432_ (.A(net3571),
    .B(_04665_),
    .C(_04824_),
    .Y(_04826_));
 sky130_fd_sc_hd__nor3_1 _22433_ (.A(_03951_),
    .B(_04825_),
    .C(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__clkinv_1 _22434_ (.A(_04824_),
    .Y(_04828_));
 sky130_fd_sc_hd__o22ai_1 _22435_ (.A1(_04651_),
    .A2(_04665_),
    .B1(_04828_),
    .B2(net3570),
    .Y(_04829_));
 sky130_fd_sc_hd__a221o_1 _22436_ (.A1(_04739_),
    .A2(_04665_),
    .B1(_04828_),
    .B2(_03951_),
    .C1(_04038_),
    .X(_04830_));
 sky130_fd_sc_hd__o21ai_0 _22437_ (.A1(net3571),
    .A2(_04829_),
    .B1(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__o21ai_0 _22438_ (.A1(_04740_),
    .A2(_04827_),
    .B1(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__xor2_1 _22439_ (.A(_03952_),
    .B(_04824_),
    .X(_04833_));
 sky130_fd_sc_hd__a22oi_2 _22440_ (.A1(_04775_),
    .A2(_04832_),
    .B1(_04833_),
    .B2(_04739_),
    .Y(_04834_));
 sky130_fd_sc_hd__nor2_2 _22441_ (.A(_04750_),
    .B(_04760_),
    .Y(_04835_));
 sky130_fd_sc_hd__maj3_1 _22442_ (.A(_04621_),
    .B(_04755_),
    .C(_04758_),
    .X(_04836_));
 sky130_fd_sc_hd__xnor2_1 _22443_ (.A(net3632),
    .B(_02856_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand2_1 _22444_ (.A(_02877_),
    .B(_03181_),
    .Y(_04838_));
 sky130_fd_sc_hd__o21ai_2 _22445_ (.A1(_02987_),
    .A2(_04837_),
    .B1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(_04751_),
    .B(_04752_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _22447_ (.A(_04751_),
    .B(_04752_),
    .Y(_04841_));
 sky130_fd_sc_hd__a21oi_2 _22448_ (.A1(_04753_),
    .A2(_04840_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__xor2_1 _22449_ (.A(_04839_),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__xnor2_1 _22450_ (.A(_04621_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__xnor2_1 _22451_ (.A(_04836_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__xnor2_1 _22452_ (.A(_04835_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__xnor2_1 _22453_ (.A(_04747_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _22454_ (.A(net3571),
    .B(_03951_),
    .Y(_04848_));
 sky130_fd_sc_hd__nor3_1 _22455_ (.A(net3628),
    .B(_04517_),
    .C(_04652_),
    .Y(_04849_));
 sky130_fd_sc_hd__o21ai_0 _22456_ (.A1(_04783_),
    .A2(_04849_),
    .B1(net3629),
    .Y(_04850_));
 sky130_fd_sc_hd__o31ai_1 _22457_ (.A1(_03470_),
    .A2(_04517_),
    .A3(_04652_),
    .B1(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21o_4 _22458_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net3668),
    .B1(net3732),
    .X(_04852_));
 sky130_fd_sc_hd__o21ai_0 _22459_ (.A1(net3627),
    .A2(_04765_),
    .B1(net3629),
    .Y(_04853_));
 sky130_fd_sc_hd__o21ai_0 _22460_ (.A1(_03460_),
    .A2(_04652_),
    .B1(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _22461_ (.A(_04652_),
    .B(_04820_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_1 _22462_ (.A(_04771_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21oi_1 _22463_ (.A1(_04852_),
    .A2(_04854_),
    .B1(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_2 _22464_ (.A(net3577),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__a31oi_4 _22465_ (.A1(net3577),
    .A2(_04781_),
    .A3(_04851_),
    .B1(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__xnor2_1 _22466_ (.A(net3570),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__nand3_1 _22467_ (.A(net3570),
    .B(_04793_),
    .C(_04859_),
    .Y(_04861_));
 sky130_fd_sc_hd__o221ai_1 _22468_ (.A1(_04848_),
    .A2(_04859_),
    .B1(_04860_),
    .B2(net3571),
    .C1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__a21oi_4 _22469_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net3668),
    .B1(net3732),
    .Y(_04863_));
 sky130_fd_sc_hd__nand3_1 _22470_ (.A(_03459_),
    .B(_03460_),
    .C(_04820_),
    .Y(_04864_));
 sky130_fd_sc_hd__o21ai_0 _22471_ (.A1(_04765_),
    .A2(_04820_),
    .B1(_03460_),
    .Y(_04865_));
 sky130_fd_sc_hd__a22o_1 _22472_ (.A1(_04852_),
    .A2(_04783_),
    .B1(_04865_),
    .B2(net3629),
    .X(_04866_));
 sky130_fd_sc_hd__nand2_1 _22473_ (.A(_04765_),
    .B(_04820_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21oi_1 _22474_ (.A1(net3628),
    .A2(_04867_),
    .B1(net3629),
    .Y(_04868_));
 sky130_fd_sc_hd__a21oi_1 _22475_ (.A1(_04820_),
    .A2(_04787_),
    .B1(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _22476_ (.A(net3577),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__o21ai_0 _22477_ (.A1(net3577),
    .A2(_04866_),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__o311ai_1 _22478_ (.A1(_03459_),
    .A2(_03460_),
    .A3(_04781_),
    .B1(_04864_),
    .C1(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__xnor2_2 _22479_ (.A(_04863_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__xnor2_1 _22480_ (.A(_04739_),
    .B(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__xnor2_1 _22481_ (.A(_04862_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__xor2_1 _22482_ (.A(_04847_),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__xnor2_1 _22483_ (.A(_04834_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__xor2_1 _22484_ (.A(_04819_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nor2_1 _22485_ (.A(_04763_),
    .B(_04795_),
    .Y(_04879_));
 sky130_fd_sc_hd__nor2_1 _22486_ (.A(_04746_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__a21oi_1 _22487_ (.A1(_04763_),
    .A2(_04795_),
    .B1(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__xnor2_1 _22488_ (.A(_04878_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21ai_2 _22489_ (.A1(_04797_),
    .A2(_04804_),
    .B1(_04805_),
    .Y(_04883_));
 sky130_fd_sc_hd__xor2_1 _22490_ (.A(_04882_),
    .B(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__o21ai_2 _22491_ (.A1(_04732_),
    .A2(_04807_),
    .B1(_04673_),
    .Y(_04885_));
 sky130_fd_sc_hd__or2_4 _22492_ (.A(_04884_),
    .B(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__nand3_1 _22493_ (.A(_04674_),
    .B(_04809_),
    .C(_04884_),
    .Y(_04887_));
 sky130_fd_sc_hd__or3_1 _22494_ (.A(_04561_),
    .B(_04598_),
    .C(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__and2_0 _22495_ (.A(net3445),
    .B(_04597_),
    .X(_04889_));
 sky130_fd_sc_hd__o21ai_0 _22496_ (.A1(_04674_),
    .A2(_04808_),
    .B1(_04809_),
    .Y(_04890_));
 sky130_fd_sc_hd__or2_0 _22497_ (.A(_04884_),
    .B(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__inv_1 _22498_ (.A(_04673_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21oi_1 _22499_ (.A1(_04892_),
    .A2(_04809_),
    .B1(_04808_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _22500_ (.A(_04884_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a21oi_1 _22501_ (.A1(_04891_),
    .A2(_04894_),
    .B1(net3670),
    .Y(_04895_));
 sky130_fd_sc_hd__o221ai_2 _22502_ (.A1(net3430),
    .A2(_04886_),
    .B1(_04888_),
    .B2(_04889_),
    .C1(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__a21oi_1 _22503_ (.A1(_02225_),
    .A2(_02942_),
    .B1(net3937),
    .Y(_04897_));
 sky130_fd_sc_hd__a22oi_2 _22504_ (.A1(net3937),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B1(_04896_),
    .B2(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__nor2_1 _22505_ (.A(net3621),
    .B(_04711_),
    .Y(_04899_));
 sky130_fd_sc_hd__nor2_1 _22506_ (.A(net3587),
    .B(_02020_),
    .Y(_04900_));
 sky130_fd_sc_hd__a211oi_1 _22507_ (.A1(net3620),
    .A2(_02020_),
    .B1(_04900_),
    .C1(net3619),
    .Y(_04901_));
 sky130_fd_sc_hd__nand2_1 _22508_ (.A(net3578),
    .B(_04686_),
    .Y(_04902_));
 sky130_fd_sc_hd__o311ai_0 _22509_ (.A1(net3578),
    .A2(_04899_),
    .A3(_04901_),
    .B1(_04902_),
    .C1(net3558),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ai_0 _22510_ (.A1(net3558),
    .A2(_03265_),
    .B1(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_1 _22511_ (.A(_02016_),
    .B(_02118_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_2 _22512_ (.A1(_02016_),
    .A2(_04904_),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__mux2i_4 _22513_ (.A0(_02953_),
    .A1(_04906_),
    .S(net3560),
    .Y(_04907_));
 sky130_fd_sc_hd__o21ai_4 _22514_ (.A1(_02171_),
    .A2(_02948_),
    .B1(_02612_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand3_1 _22515_ (.A(net3726),
    .B(_10393_),
    .C(net3587),
    .Y(_04909_));
 sky130_fd_sc_hd__o21ai_0 _22516_ (.A1(net3587),
    .A2(_03272_),
    .B1(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__a21oi_1 _22517_ (.A1(net3587),
    .A2(_03272_),
    .B1(_10393_),
    .Y(_04911_));
 sky130_fd_sc_hd__a21oi_1 _22518_ (.A1(_02127_),
    .A2(_04910_),
    .B1(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__a221oi_1 _22519_ (.A1(net3603),
    .A2(_04907_),
    .B1(_04908_),
    .B2(net3602),
    .C1(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__o21ai_2 _22520_ (.A1(net3471),
    .A2(_02702_),
    .B1(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_4 _22521_ (.A(net3744),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__o2111ai_2 _22522_ (.A1(net321),
    .A2(net3415),
    .B1(_04915_),
    .C1(_11563_),
    .D1(net3469),
    .Y(_04916_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_381 ();
 sky130_fd_sc_hd__nand2_1 _22524_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_02842_),
    .Y(_04918_));
 sky130_fd_sc_hd__o21ai_2 _22525_ (.A1(net3822),
    .A2(_02841_),
    .B1(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21oi_4 _22526_ (.A1(_01670_),
    .A2(_04919_),
    .B1(_03289_),
    .Y(_04920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_380 ();
 sky130_fd_sc_hd__nor2_1 _22528_ (.A(_02153_),
    .B(_04920_),
    .Y(_04922_));
 sky130_fd_sc_hd__a22o_1 _22529_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .A2(_02153_),
    .B1(net3403),
    .B2(_04922_),
    .X(_00539_));
 sky130_fd_sc_hd__nand3_1 _22530_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_02419_),
    .C(net41),
    .Y(_04923_));
 sky130_fd_sc_hd__nand3_1 _22531_ (.A(_02423_),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .C(net32),
    .Y(_04924_));
 sky130_fd_sc_hd__a221oi_1 _22532_ (.A1(\load_store_unit_i.rdata_q[14] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[6] ),
    .C1(_02847_),
    .Y(_04925_));
 sky130_fd_sc_hd__a31oi_1 _22533_ (.A1(_02847_),
    .A2(_04923_),
    .A3(_04924_),
    .B1(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__and3_1 _22534_ (.A(_02423_),
    .B(_02419_),
    .C(net55),
    .X(_04927_));
 sky130_fd_sc_hd__a22oi_1 _22535_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net50),
    .B1(_03238_),
    .B2(\load_store_unit_i.rdata_q[22] ),
    .Y(_04928_));
 sky130_fd_sc_hd__nor2_1 _22536_ (.A(_03237_),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__a22oi_1 _22537_ (.A1(net3602),
    .A2(_04231_),
    .B1(_04233_),
    .B2(net3603),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _22538_ (.A(_08000_),
    .B(_02127_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_1 _22539_ (.A(net3601),
    .B(_02129_),
    .Y(_04932_));
 sky130_fd_sc_hd__o21ai_0 _22540_ (.A1(net3601),
    .A2(_02136_),
    .B1(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__a32oi_2 _22541_ (.A1(net3601),
    .A2(_03272_),
    .A3(_04931_),
    .B1(_04933_),
    .B2(_08000_),
    .Y(_04934_));
 sky130_fd_sc_hd__o211ai_1 _22542_ (.A1(net3529),
    .A2(_02702_),
    .B1(_04930_),
    .C1(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__mux2i_2 _22543_ (.A0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A1(_03885_),
    .S(_02000_),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_1 _22544_ (.A(net3937),
    .B(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .Y(_04937_));
 sky130_fd_sc_hd__o211ai_1 _22545_ (.A1(net3937),
    .A2(_04936_),
    .B1(_04937_),
    .C1(_07857_),
    .Y(_04938_));
 sky130_fd_sc_hd__o21ai_4 _22546_ (.A1(net3739),
    .A2(_04935_),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand3_4 _22547_ (.A(_11662_),
    .B(_01655_),
    .C(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__o41ai_2 _22548_ (.A1(net3469),
    .A2(_04926_),
    .A3(_04927_),
    .A4(_04929_),
    .B1(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_379 ();
 sky130_fd_sc_hd__nand2_1 _22550_ (.A(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .B(_03280_),
    .Y(_04943_));
 sky130_fd_sc_hd__o21ai_0 _22551_ (.A1(_03280_),
    .A2(net3444),
    .B1(_04943_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _22552_ (.A(net3530),
    .B(_02006_),
    .Y(_04944_));
 sky130_fd_sc_hd__mux2i_1 _22553_ (.A0(_02136_),
    .A1(_02133_),
    .S(_08810_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _22554_ (.A(_08810_),
    .B(_03272_),
    .Y(_04946_));
 sky130_fd_sc_hd__a21oi_1 _22555_ (.A1(_08779_),
    .A2(_02127_),
    .B1(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__a221oi_1 _22556_ (.A1(net3602),
    .A2(_04112_),
    .B1(_04945_),
    .B2(_08779_),
    .C1(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__o211ai_1 _22557_ (.A1(_02020_),
    .A2(_04106_),
    .B1(_04944_),
    .C1(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand2_1 _22558_ (.A(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B(_02225_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _22559_ (.A(_02000_),
    .B(_03903_),
    .Y(_04951_));
 sky130_fd_sc_hd__nand2_2 _22560_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__mux2i_1 _22561_ (.A0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A1(_04952_),
    .S(_08009_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand2_4 _22562_ (.A(net3756),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__o21ai_2 _22563_ (.A1(_08316_),
    .A2(_04949_),
    .B1(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__and3_1 _22564_ (.A(_02423_),
    .B(\load_store_unit_i.rdata_offset_q[0] ),
    .C(net33),
    .X(_04956_));
 sky130_fd_sc_hd__a21oi_1 _22565_ (.A1(net42),
    .A2(_02424_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__a221oi_1 _22566_ (.A1(\load_store_unit_i.rdata_q[15] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[7] ),
    .C1(_02847_),
    .Y(_04958_));
 sky130_fd_sc_hd__a21oi_1 _22567_ (.A1(_02847_),
    .A2(_04957_),
    .B1(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nor2_4 _22568_ (.A(_10666_),
    .B(_03237_),
    .Y(_04960_));
 sky130_fd_sc_hd__nor2_4 _22569_ (.A(_02417_),
    .B(_03237_),
    .Y(_04961_));
 sky130_fd_sc_hd__a22o_1 _22570_ (.A1(net51),
    .A2(_04960_),
    .B1(_04961_),
    .B2(\load_store_unit_i.rdata_q[23] ),
    .X(_04962_));
 sky130_fd_sc_hd__a2111oi_1 _22571_ (.A1(net56),
    .A2(_02418_),
    .B1(_04959_),
    .C1(_04962_),
    .D1(net3469),
    .Y(_04963_));
 sky130_fd_sc_hd__a31o_4 _22572_ (.A1(_11683_),
    .A2(net3469),
    .A3(_04955_),
    .B1(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_378 ();
 sky130_fd_sc_hd__nand2_1 _22574_ (.A(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .B(_03280_),
    .Y(_04966_));
 sky130_fd_sc_hd__o21ai_0 _22575_ (.A1(_03280_),
    .A2(_04964_),
    .B1(_04966_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _22576_ (.A(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .B(_03280_),
    .Y(_04967_));
 sky130_fd_sc_hd__o21ai_0 _22577_ (.A1(_02145_),
    .A2(_03280_),
    .B1(_04967_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _22578_ (.A(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .B(_03280_),
    .Y(_04968_));
 sky130_fd_sc_hd__o21ai_0 _22579_ (.A1(_02297_),
    .A2(_03280_),
    .B1(_04968_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _22580_ (.A(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .B(_03280_),
    .Y(_04969_));
 sky130_fd_sc_hd__o21ai_0 _22581_ (.A1(_02414_),
    .A2(_03280_),
    .B1(_04969_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _22582_ (.A(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .B(_03280_),
    .Y(_04970_));
 sky130_fd_sc_hd__o21ai_0 _22583_ (.A1(_02535_),
    .A2(_03280_),
    .B1(_04970_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _22584_ (.A(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .B(_03280_),
    .Y(_04971_));
 sky130_fd_sc_hd__o21ai_0 _22585_ (.A1(_02628_),
    .A2(_03280_),
    .B1(_04971_),
    .Y(_00546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_377 ();
 sky130_fd_sc_hd__nand2_1 _22587_ (.A(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .B(_03280_),
    .Y(_04973_));
 sky130_fd_sc_hd__o21ai_0 _22588_ (.A1(net3453),
    .A2(_03280_),
    .B1(_04973_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _22589_ (.A(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .B(_03280_),
    .Y(_04974_));
 sky130_fd_sc_hd__o21ai_0 _22590_ (.A1(_02837_),
    .A2(_03280_),
    .B1(_04974_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _22591_ (.A(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .B(_03280_),
    .Y(_04975_));
 sky130_fd_sc_hd__o21ai_0 _22592_ (.A1(_02963_),
    .A2(_03280_),
    .B1(_04975_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _22593_ (.A(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .B(_03280_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_0 _22594_ (.A1(net3447),
    .A2(_03280_),
    .B1(_04976_),
    .Y(_00550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_376 ();
 sky130_fd_sc_hd__or3_4 _22596_ (.A(net3946),
    .B(net3827),
    .C(net3945),
    .X(_04978_));
 sky130_fd_sc_hd__nor2_4 _22597_ (.A(_04978_),
    .B(_03094_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _22598_ (.A(net3446),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _22599_ (.A(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .B(_03280_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _22600_ (.A(_04980_),
    .B(_04981_),
    .Y(_00551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_375 ();
 sky130_fd_sc_hd__nand2_1 _22602_ (.A(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .B(_03280_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ai_0 _22603_ (.A1(_03280_),
    .A2(net3425),
    .B1(_04983_),
    .Y(_00552_));
 sky130_fd_sc_hd__mux2_1 _22604_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .A1(net3416),
    .S(_04979_),
    .X(_00553_));
 sky130_fd_sc_hd__nand2_1 _22605_ (.A(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .B(_03280_),
    .Y(_04984_));
 sky130_fd_sc_hd__o21ai_0 _22606_ (.A1(_03280_),
    .A2(net3433),
    .B1(_04984_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _22607_ (.A(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .B(_03280_),
    .Y(_04985_));
 sky130_fd_sc_hd__o21ai_0 _22608_ (.A1(_03280_),
    .A2(net3413),
    .B1(_04985_),
    .Y(_00555_));
 sky130_fd_sc_hd__mux2_1 _22609_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .A1(net3412),
    .S(_04979_),
    .X(_00556_));
 sky130_fd_sc_hd__nand2_1 _22610_ (.A(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .B(_03280_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_0 _22611_ (.A1(_03280_),
    .A2(net3411),
    .B1(_04986_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _22612_ (.A(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .B(_03280_),
    .Y(_04987_));
 sky130_fd_sc_hd__o21ai_0 _22613_ (.A1(_03280_),
    .A2(net3410),
    .B1(_04987_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _22614_ (.A(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .B(_03280_),
    .Y(_04988_));
 sky130_fd_sc_hd__o21ai_0 _22615_ (.A1(_03280_),
    .A2(net3409),
    .B1(_04988_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _22616_ (.A(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .B(_03280_),
    .Y(_04989_));
 sky130_fd_sc_hd__o21ai_0 _22617_ (.A1(_03280_),
    .A2(net3408),
    .B1(_04989_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _22618_ (.A(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .B(_03280_),
    .Y(_04990_));
 sky130_fd_sc_hd__o21ai_0 _22619_ (.A1(_03280_),
    .A2(net3407),
    .B1(_04990_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _22620_ (.A(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .B(_03280_),
    .Y(_04991_));
 sky130_fd_sc_hd__o21ai_0 _22621_ (.A1(_03280_),
    .A2(net3406),
    .B1(_04991_),
    .Y(_00562_));
 sky130_fd_sc_hd__nor2_1 _22622_ (.A(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .B(_04979_),
    .Y(_04992_));
 sky130_fd_sc_hd__a31oi_1 _22623_ (.A1(_04979_),
    .A2(net3405),
    .A3(net3457),
    .B1(_04992_),
    .Y(_00563_));
 sky130_fd_sc_hd__mux2_1 _22624_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .A1(net3404),
    .S(_04979_),
    .X(_00564_));
 sky130_fd_sc_hd__nor2_1 _22625_ (.A(_03280_),
    .B(_04920_),
    .Y(_04993_));
 sky130_fd_sc_hd__a22o_1 _22626_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .A2(_03280_),
    .B1(net3403),
    .B2(_04993_),
    .X(_00565_));
 sky130_fd_sc_hd__a22oi_1 _22627_ (.A1(\load_store_unit_i.rdata_q[8] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[0] ),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_1 _22628_ (.A(_02419_),
    .B(net34),
    .Y(_04995_));
 sky130_fd_sc_hd__a21oi_1 _22629_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net57),
    .B1(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_04996_));
 sky130_fd_sc_hd__a21oi_1 _22630_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_04995_),
    .B1(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a222oi_1 _22631_ (.A1(net27),
    .A2(_02418_),
    .B1(_04960_),
    .B2(net43),
    .C1(_04997_),
    .C2(_02847_),
    .Y(_04998_));
 sky130_fd_sc_hd__nand2_1 _22632_ (.A(\load_store_unit_i.rdata_q[16] ),
    .B(_04961_),
    .Y(_04999_));
 sky130_fd_sc_hd__o2111ai_4 _22633_ (.A1(_02847_),
    .A2(_04994_),
    .B1(_04998_),
    .C1(_04999_),
    .D1(net3472),
    .Y(_05000_));
 sky130_fd_sc_hd__nor2b_2 _22634_ (.A(_04470_),
    .B_N(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .Y(_05001_));
 sky130_fd_sc_hd__a211oi_4 _22635_ (.A1(_02977_),
    .A2(_04470_),
    .B1(_05001_),
    .C1(_08498_),
    .Y(_05002_));
 sky130_fd_sc_hd__nand2_4 _22636_ (.A(net3462),
    .B(net3461),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _22637_ (.A(net3603),
    .B(_04908_),
    .Y(_05004_));
 sky130_fd_sc_hd__xor2_1 _22638_ (.A(net3596),
    .B(_02133_),
    .X(_05005_));
 sky130_fd_sc_hd__a21oi_1 _22639_ (.A1(net3621),
    .A2(net3620),
    .B1(_03273_),
    .Y(_05006_));
 sky130_fd_sc_hd__o21ai_0 _22640_ (.A1(_02184_),
    .A2(_05005_),
    .B1(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__o2111ai_2 _22641_ (.A1(_10701_),
    .A2(_02702_),
    .B1(_05004_),
    .C1(_05007_),
    .D1(net3737),
    .Y(_05008_));
 sky130_fd_sc_hd__a221oi_4 _22642_ (.A1(net372),
    .A2(_05003_),
    .B1(net3602),
    .B2(_04907_),
    .C1(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__o311ai_4 _22643_ (.A1(net3738),
    .A2(_05002_),
    .A3(_05009_),
    .B1(_11040_),
    .C1(net3469),
    .Y(_05010_));
 sky130_fd_sc_hd__nand2_8 _22644_ (.A(_05000_),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_374 ();
 sky130_fd_sc_hd__nor3b_4 _22646_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .C_N(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Y(_05013_));
 sky130_fd_sc_hd__nor2b_4 _22647_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .B_N(_02150_),
    .Y(_05014_));
 sky130_fd_sc_hd__nor2b_4 _22648_ (.A(net3828),
    .B_N(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_8 _22649_ (.A(_05013_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_371 ();
 sky130_fd_sc_hd__nand2_1 _22653_ (.A(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .B(_05016_),
    .Y(_05020_));
 sky130_fd_sc_hd__o21ai_0 _22654_ (.A1(_05011_),
    .A2(_05016_),
    .B1(_05020_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _22655_ (.A(net3597),
    .B(net308),
    .Y(_05021_));
 sky130_fd_sc_hd__xnor2_1 _22656_ (.A(_02133_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__o221ai_1 _22657_ (.A1(net3597),
    .A2(net308),
    .B1(_02184_),
    .B2(_05022_),
    .C1(_02137_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21ai_0 _22658_ (.A1(_13118_),
    .A2(_02702_),
    .B1(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__a221oi_1 _22659_ (.A1(net3602),
    .A2(_04716_),
    .B1(_04717_),
    .B2(net3603),
    .C1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_1 _22660_ (.A(net3746),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _22661_ (.A(_03104_),
    .B(_04470_),
    .Y(_05027_));
 sky130_fd_sc_hd__o21ai_4 _22662_ (.A1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A2(_04470_),
    .B1(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__nand2_2 _22663_ (.A(net3739),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__a21oi_2 _22664_ (.A1(_05026_),
    .A2(_05029_),
    .B1(net3738),
    .Y(_05030_));
 sky130_fd_sc_hd__a21oi_4 _22665_ (.A1(net3738),
    .A2(_11352_),
    .B1(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__a22oi_1 _22666_ (.A1(\load_store_unit_i.rdata_q[9] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[1] ),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _22667_ (.A(_02419_),
    .B(net35),
    .Y(_05033_));
 sky130_fd_sc_hd__a21oi_1 _22668_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net58),
    .B1(net3822),
    .Y(_05034_));
 sky130_fd_sc_hd__a21oi_1 _22669_ (.A1(net3822),
    .A2(_05033_),
    .B1(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__a222oi_1 _22670_ (.A1(net38),
    .A2(_02418_),
    .B1(_04960_),
    .B2(net44),
    .C1(_05035_),
    .C2(_02847_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _22671_ (.A(\load_store_unit_i.rdata_q[17] ),
    .B(_04961_),
    .Y(_05037_));
 sky130_fd_sc_hd__o2111ai_2 _22672_ (.A1(_02847_),
    .A2(_05032_),
    .B1(_05036_),
    .C1(_05037_),
    .D1(net3472),
    .Y(_05038_));
 sky130_fd_sc_hd__o21ai_4 _22673_ (.A1(net3472),
    .A2(_05031_),
    .B1(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_370 ();
 sky130_fd_sc_hd__nand2_1 _22675_ (.A(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .B(_05016_),
    .Y(_05041_));
 sky130_fd_sc_hd__o21ai_0 _22676_ (.A1(_05016_),
    .A2(_05039_),
    .B1(_05041_),
    .Y(_00567_));
 sky130_fd_sc_hd__a22oi_1 _22677_ (.A1(\load_store_unit_i.rdata_q[10] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[2] ),
    .Y(_05042_));
 sky130_fd_sc_hd__nor2_1 _22678_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_03286_),
    .Y(_05043_));
 sky130_fd_sc_hd__a21oi_1 _22679_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03284_),
    .B1(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__a222oi_1 _22680_ (.A1(net49),
    .A2(_02418_),
    .B1(_04960_),
    .B2(net45),
    .C1(_05044_),
    .C2(_02847_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _22681_ (.A(\load_store_unit_i.rdata_q[18] ),
    .B(_04961_),
    .Y(_05046_));
 sky130_fd_sc_hd__o2111ai_4 _22682_ (.A1(_02847_),
    .A2(_05042_),
    .B1(_05045_),
    .C1(_05046_),
    .D1(net3472),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _22683_ (.A(net3598),
    .B(net3622),
    .Y(_05048_));
 sky130_fd_sc_hd__nor2_1 _22684_ (.A(net3598),
    .B(net3622),
    .Y(_05049_));
 sky130_fd_sc_hd__xnor2_1 _22685_ (.A(_05049_),
    .B(_02133_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2_1 _22686_ (.A(_02127_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__a32o_1 _22687_ (.A1(_05048_),
    .A2(_02137_),
    .A3(_05051_),
    .B1(_04693_),
    .B2(net3603),
    .X(_05052_));
 sky130_fd_sc_hd__a221o_4 _22688_ (.A1(net171),
    .A2(_02006_),
    .B1(net3602),
    .B2(_04692_),
    .C1(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o21ai_1 _22689_ (.A1(net3937),
    .A2(_02225_),
    .B1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_2 _22690_ (.A(_03401_),
    .B(_04470_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand3_4 _22691_ (.A(net3756),
    .B(_05054_),
    .C(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__o21ai_2 _22692_ (.A1(net3739),
    .A2(_05053_),
    .B1(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand3_4 _22693_ (.A(_11080_),
    .B(_01655_),
    .C(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_8 _22694_ (.A(_05047_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_369 ();
 sky130_fd_sc_hd__nand2_1 _22696_ (.A(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .B(_05016_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21ai_0 _22697_ (.A1(_05016_),
    .A2(_05059_),
    .B1(_05061_),
    .Y(_00568_));
 sky130_fd_sc_hd__nor2_1 _22698_ (.A(net3623),
    .B(net3599),
    .Y(_05062_));
 sky130_fd_sc_hd__xor2_1 _22699_ (.A(_02133_),
    .B(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__nand2_1 _22700_ (.A(net3623),
    .B(net3599),
    .Y(_05064_));
 sky130_fd_sc_hd__o211ai_1 _22701_ (.A1(_02184_),
    .A2(_05063_),
    .B1(_05064_),
    .C1(_02137_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21ai_2 _22702_ (.A1(net3534),
    .A2(_02702_),
    .B1(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__a221oi_4 _22703_ (.A1(net3602),
    .A2(_04581_),
    .B1(_04585_),
    .B2(net3603),
    .C1(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_2 _22704_ (.A(_02000_),
    .B(_03418_),
    .Y(_05068_));
 sky130_fd_sc_hd__o21ai_2 _22705_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_02000_),
    .B1(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__nor2_4 _22706_ (.A(net3937),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__a211oi_2 _22707_ (.A1(net3937),
    .A2(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B1(net3748),
    .C1(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__a21oi_2 _22708_ (.A1(_08498_),
    .A2(_05067_),
    .B1(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__a22oi_1 _22709_ (.A1(\load_store_unit_i.rdata_q[11] ),
    .A2(_02424_),
    .B1(_02420_),
    .B2(\load_store_unit_i.rdata_q[3] ),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _22710_ (.A(_02419_),
    .B(net37),
    .Y(_05074_));
 sky130_fd_sc_hd__a21oi_1 _22711_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net29),
    .B1(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_05075_));
 sky130_fd_sc_hd__a21oi_1 _22712_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_05074_),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a222oi_1 _22713_ (.A1(net52),
    .A2(_02418_),
    .B1(_05076_),
    .B2(_02847_),
    .C1(_04961_),
    .C2(\load_store_unit_i.rdata_q[19] ),
    .Y(_05077_));
 sky130_fd_sc_hd__nand2_1 _22714_ (.A(net46),
    .B(_04960_),
    .Y(_05078_));
 sky130_fd_sc_hd__o2111ai_1 _22715_ (.A1(_02847_),
    .A2(_05073_),
    .B1(_05077_),
    .C1(_05078_),
    .D1(net3472),
    .Y(_05079_));
 sky130_fd_sc_hd__o31ai_2 _22716_ (.A1(_11610_),
    .A2(net3472),
    .A3(_05072_),
    .B1(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_368 ();
 sky130_fd_sc_hd__nand2_1 _22718_ (.A(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .B(_05016_),
    .Y(_05082_));
 sky130_fd_sc_hd__o21ai_0 _22719_ (.A1(_05016_),
    .A2(net3463),
    .B1(_05082_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _22720_ (.A(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .B(_05016_),
    .Y(_05083_));
 sky130_fd_sc_hd__o21ai_0 _22721_ (.A1(net3459),
    .A2(_05016_),
    .B1(_05083_),
    .Y(_00570_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_367 ();
 sky130_fd_sc_hd__nand2_1 _22723_ (.A(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .B(_05016_),
    .Y(_05085_));
 sky130_fd_sc_hd__o21ai_0 _22724_ (.A1(_04483_),
    .A2(_05016_),
    .B1(_05085_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _22725_ (.A(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .B(_05016_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_0 _22726_ (.A1(net3444),
    .A2(_05016_),
    .B1(_05086_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _22727_ (.A(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .B(_05016_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21ai_0 _22728_ (.A1(_04964_),
    .A2(_05016_),
    .B1(_05087_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _22729_ (.A(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .B(_05016_),
    .Y(_05088_));
 sky130_fd_sc_hd__o21ai_0 _22730_ (.A1(_02145_),
    .A2(_05016_),
    .B1(_05088_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _22731_ (.A(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .B(_05016_),
    .Y(_05089_));
 sky130_fd_sc_hd__o21ai_0 _22732_ (.A1(_02297_),
    .A2(_05016_),
    .B1(_05089_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _22733_ (.A(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .B(_05016_),
    .Y(_05090_));
 sky130_fd_sc_hd__o21ai_0 _22734_ (.A1(_02414_),
    .A2(_05016_),
    .B1(_05090_),
    .Y(_00576_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_366 ();
 sky130_fd_sc_hd__nand2_1 _22736_ (.A(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .B(_05016_),
    .Y(_05092_));
 sky130_fd_sc_hd__o21ai_0 _22737_ (.A1(_02535_),
    .A2(_05016_),
    .B1(_05092_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _22738_ (.A(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .B(_05016_),
    .Y(_05093_));
 sky130_fd_sc_hd__o21ai_0 _22739_ (.A1(_02628_),
    .A2(_05016_),
    .B1(_05093_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _22740_ (.A(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .B(_05016_),
    .Y(_05094_));
 sky130_fd_sc_hd__o21ai_0 _22741_ (.A1(net3453),
    .A2(_05016_),
    .B1(_05094_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _22742_ (.A(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .B(_05016_),
    .Y(_05095_));
 sky130_fd_sc_hd__o21ai_0 _22743_ (.A1(_02837_),
    .A2(_05016_),
    .B1(_05095_),
    .Y(_00580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_365 ();
 sky130_fd_sc_hd__nand2_1 _22745_ (.A(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .B(_05016_),
    .Y(_05097_));
 sky130_fd_sc_hd__o21ai_0 _22746_ (.A1(_02963_),
    .A2(_05016_),
    .B1(_05097_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _22747_ (.A(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .B(_05016_),
    .Y(_05098_));
 sky130_fd_sc_hd__o21ai_0 _22748_ (.A1(net3447),
    .A2(_05016_),
    .B1(_05098_),
    .Y(_00582_));
 sky130_fd_sc_hd__or3b_4 _22749_ (.A(net3946),
    .B(net3945),
    .C_N(net3827),
    .X(_05099_));
 sky130_fd_sc_hd__nand2b_4 _22750_ (.A_N(net3828),
    .B(_05014_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_4 _22751_ (.A(_05099_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand2_1 _22752_ (.A(net3446),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _22753_ (.A(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .B(_05016_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _22754_ (.A(_05102_),
    .B(_05103_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _22755_ (.A(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .B(_05016_),
    .Y(_05104_));
 sky130_fd_sc_hd__o21ai_0 _22756_ (.A1(net3425),
    .A2(_05016_),
    .B1(_05104_),
    .Y(_00584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_364 ();
 sky130_fd_sc_hd__nand2_1 _22758_ (.A(net3416),
    .B(_05101_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_1 _22759_ (.A(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .B(_05016_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand2_1 _22760_ (.A(_05106_),
    .B(_05107_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _22761_ (.A(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .B(_05016_),
    .Y(_05108_));
 sky130_fd_sc_hd__o21ai_0 _22762_ (.A1(net3433),
    .A2(_05016_),
    .B1(_05108_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _22763_ (.A(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .B(_05016_),
    .Y(_05109_));
 sky130_fd_sc_hd__o21ai_0 _22764_ (.A1(net3413),
    .A2(_05016_),
    .B1(_05109_),
    .Y(_00587_));
 sky130_fd_sc_hd__mux2_1 _22765_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A1(net3412),
    .S(_05101_),
    .X(_00588_));
 sky130_fd_sc_hd__nand2_1 _22766_ (.A(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .B(_05016_),
    .Y(_05110_));
 sky130_fd_sc_hd__o21ai_0 _22767_ (.A1(net3411),
    .A2(_05016_),
    .B1(_05110_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .B(_05016_),
    .Y(_05111_));
 sky130_fd_sc_hd__o21ai_0 _22769_ (.A1(net3410),
    .A2(_05016_),
    .B1(_05111_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _22770_ (.A(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .B(_05016_),
    .Y(_05112_));
 sky130_fd_sc_hd__o21ai_0 _22771_ (.A1(net3409),
    .A2(_05016_),
    .B1(_05112_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _22772_ (.A(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .B(_05016_),
    .Y(_05113_));
 sky130_fd_sc_hd__o21ai_0 _22773_ (.A1(net3408),
    .A2(_05016_),
    .B1(_05113_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _22774_ (.A(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .B(_05016_),
    .Y(_05114_));
 sky130_fd_sc_hd__o21ai_0 _22775_ (.A1(net3407),
    .A2(_05016_),
    .B1(_05114_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _22776_ (.A(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .B(_05016_),
    .Y(_05115_));
 sky130_fd_sc_hd__o21ai_0 _22777_ (.A1(net3406),
    .A2(_05016_),
    .B1(_05115_),
    .Y(_00594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_362 ();
 sky130_fd_sc_hd__nor2_1 _22780_ (.A(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .B(_05101_),
    .Y(_05118_));
 sky130_fd_sc_hd__a31oi_1 _22781_ (.A1(net3405),
    .A2(net3457),
    .A3(_05101_),
    .B1(_05118_),
    .Y(_00595_));
 sky130_fd_sc_hd__mux2_1 _22782_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(net3404),
    .S(_05101_),
    .X(_00596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_361 ();
 sky130_fd_sc_hd__nor2_1 _22784_ (.A(_04920_),
    .B(_05016_),
    .Y(_05120_));
 sky130_fd_sc_hd__a22o_1 _22785_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A2(_05016_),
    .B1(_05120_),
    .B2(net3403),
    .X(_00597_));
 sky130_fd_sc_hd__nand2_2 _22786_ (.A(net3829),
    .B(_02150_),
    .Y(_05121_));
 sky130_fd_sc_hd__nor2_4 _22787_ (.A(net3828),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_8 _22788_ (.A(_05013_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_358 ();
 sky130_fd_sc_hd__nand2_1 _22792_ (.A(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .B(_05123_),
    .Y(_05127_));
 sky130_fd_sc_hd__o21ai_0 _22793_ (.A1(_05011_),
    .A2(_05123_),
    .B1(_05127_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _22794_ (.A(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .B(_05123_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_0 _22795_ (.A1(_05039_),
    .A2(_05123_),
    .B1(_05128_),
    .Y(_00599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_357 ();
 sky130_fd_sc_hd__nand2_1 _22797_ (.A(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .B(_05123_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_0 _22798_ (.A1(_05059_),
    .A2(_05123_),
    .B1(_05130_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _22799_ (.A(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .B(_05123_),
    .Y(_05131_));
 sky130_fd_sc_hd__o21ai_0 _22800_ (.A1(net3463),
    .A2(_05123_),
    .B1(_05131_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _22801_ (.A(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .B(_05123_),
    .Y(_05132_));
 sky130_fd_sc_hd__o21ai_0 _22802_ (.A1(net3459),
    .A2(_05123_),
    .B1(_05132_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _22803_ (.A(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .B(_05123_),
    .Y(_05133_));
 sky130_fd_sc_hd__o21ai_0 _22804_ (.A1(_04483_),
    .A2(_05123_),
    .B1(_05133_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _22805_ (.A(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .B(_05123_),
    .Y(_05134_));
 sky130_fd_sc_hd__o21ai_0 _22806_ (.A1(net3444),
    .A2(_05123_),
    .B1(_05134_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _22807_ (.A(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .B(_05123_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_0 _22808_ (.A1(_04964_),
    .A2(_05123_),
    .B1(_05135_),
    .Y(_00605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_356 ();
 sky130_fd_sc_hd__nand2_1 _22810_ (.A(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .B(_05123_),
    .Y(_05137_));
 sky130_fd_sc_hd__o21ai_0 _22811_ (.A1(_02145_),
    .A2(_05123_),
    .B1(_05137_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _22812_ (.A(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .B(_05123_),
    .Y(_05138_));
 sky130_fd_sc_hd__o21ai_0 _22813_ (.A1(_02297_),
    .A2(_05123_),
    .B1(_05138_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .B(_05123_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_0 _22815_ (.A1(_02414_),
    .A2(_05123_),
    .B1(_05139_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _22816_ (.A(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .B(_05123_),
    .Y(_05140_));
 sky130_fd_sc_hd__o21ai_0 _22817_ (.A1(_02535_),
    .A2(_05123_),
    .B1(_05140_),
    .Y(_00609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_355 ();
 sky130_fd_sc_hd__nand2_1 _22819_ (.A(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .B(_05123_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_0 _22820_ (.A1(_02628_),
    .A2(_05123_),
    .B1(_05142_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _22821_ (.A(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .B(_05123_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21ai_0 _22822_ (.A1(net3453),
    .A2(_05123_),
    .B1(_05143_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _22823_ (.A(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .B(_05123_),
    .Y(_05144_));
 sky130_fd_sc_hd__o21ai_0 _22824_ (.A1(_02837_),
    .A2(_05123_),
    .B1(_05144_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _22825_ (.A(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .B(_05123_),
    .Y(_05145_));
 sky130_fd_sc_hd__o21ai_0 _22826_ (.A1(_02963_),
    .A2(_05123_),
    .B1(_05145_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _22827_ (.A(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .B(_05123_),
    .Y(_05146_));
 sky130_fd_sc_hd__o21ai_0 _22828_ (.A1(net3447),
    .A2(_05123_),
    .B1(_05146_),
    .Y(_00614_));
 sky130_fd_sc_hd__or2_4 _22829_ (.A(net3828),
    .B(_05121_),
    .X(_05147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_354 ();
 sky130_fd_sc_hd__nor2_4 _22831_ (.A(_05099_),
    .B(_05147_),
    .Y(_05149_));
 sky130_fd_sc_hd__nand2_1 _22832_ (.A(net3446),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_1 _22833_ (.A(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .B(_05123_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _22834_ (.A(_05150_),
    .B(_05151_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _22835_ (.A(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .B(_05123_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_0 _22836_ (.A1(net3425),
    .A2(_05123_),
    .B1(_05152_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _22837_ (.A(net3416),
    .B(_05149_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand2_1 _22838_ (.A(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .B(_05123_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(_05153_),
    .B(_05154_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _22840_ (.A(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .B(_05123_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21ai_0 _22841_ (.A1(net3433),
    .A2(_05123_),
    .B1(_05155_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _22842_ (.A(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .B(_05123_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_0 _22843_ (.A1(net3413),
    .A2(_05123_),
    .B1(_05156_),
    .Y(_00619_));
 sky130_fd_sc_hd__mux2_1 _22844_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A1(net3412),
    .S(_05149_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _22845_ (.A(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .B(_05123_),
    .Y(_05157_));
 sky130_fd_sc_hd__o21ai_0 _22846_ (.A1(net3411),
    .A2(_05123_),
    .B1(_05157_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _22847_ (.A(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .B(_05123_),
    .Y(_05158_));
 sky130_fd_sc_hd__o21ai_0 _22848_ (.A1(net3410),
    .A2(_05123_),
    .B1(_05158_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _22849_ (.A(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .B(_05123_),
    .Y(_05159_));
 sky130_fd_sc_hd__o21ai_0 _22850_ (.A1(net3409),
    .A2(_05123_),
    .B1(_05159_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _22851_ (.A(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .B(_05123_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21ai_0 _22852_ (.A1(net3408),
    .A2(_05123_),
    .B1(_05160_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _22853_ (.A(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .B(_05123_),
    .Y(_05161_));
 sky130_fd_sc_hd__o21ai_0 _22854_ (.A1(net3407),
    .A2(_05123_),
    .B1(_05161_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _22855_ (.A(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .B(_05123_),
    .Y(_05162_));
 sky130_fd_sc_hd__o21ai_0 _22856_ (.A1(net3406),
    .A2(_05123_),
    .B1(_05162_),
    .Y(_00626_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .B(_05149_),
    .Y(_05163_));
 sky130_fd_sc_hd__a31oi_1 _22858_ (.A1(net3405),
    .A2(net3457),
    .A3(_05149_),
    .B1(_05163_),
    .Y(_00627_));
 sky130_fd_sc_hd__mux2_1 _22859_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A1(net3404),
    .S(_05149_),
    .X(_00628_));
 sky130_fd_sc_hd__nor2_1 _22860_ (.A(_04920_),
    .B(_05123_),
    .Y(_05164_));
 sky130_fd_sc_hd__a22o_1 _22861_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(_05123_),
    .B1(_05164_),
    .B2(net3403),
    .X(_00629_));
 sky130_fd_sc_hd__and2_4 _22862_ (.A(net3828),
    .B(_05014_),
    .X(_05165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_353 ();
 sky130_fd_sc_hd__nand2_8 _22864_ (.A(_05013_),
    .B(_05165_),
    .Y(_05167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_350 ();
 sky130_fd_sc_hd__nand2_1 _22868_ (.A(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .B(_05167_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_0 _22869_ (.A1(_05011_),
    .A2(_05167_),
    .B1(_05171_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _22870_ (.A(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .B(_05167_),
    .Y(_05172_));
 sky130_fd_sc_hd__o21ai_0 _22871_ (.A1(_05039_),
    .A2(_05167_),
    .B1(_05172_),
    .Y(_00631_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_349 ();
 sky130_fd_sc_hd__nand2_1 _22873_ (.A(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .B(_05167_),
    .Y(_05174_));
 sky130_fd_sc_hd__o21ai_0 _22874_ (.A1(_05059_),
    .A2(_05167_),
    .B1(_05174_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _22875_ (.A(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .B(_05167_),
    .Y(_05175_));
 sky130_fd_sc_hd__o21ai_0 _22876_ (.A1(net3463),
    .A2(_05167_),
    .B1(_05175_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _22877_ (.A(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .B(_05167_),
    .Y(_05176_));
 sky130_fd_sc_hd__o21ai_0 _22878_ (.A1(net3459),
    .A2(_05167_),
    .B1(_05176_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _22879_ (.A(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .B(_05167_),
    .Y(_05177_));
 sky130_fd_sc_hd__o21ai_0 _22880_ (.A1(_04483_),
    .A2(_05167_),
    .B1(_05177_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _22881_ (.A(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .B(_05167_),
    .Y(_05178_));
 sky130_fd_sc_hd__o21ai_0 _22882_ (.A1(net3444),
    .A2(_05167_),
    .B1(_05178_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _22883_ (.A(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .B(_05167_),
    .Y(_05179_));
 sky130_fd_sc_hd__o21ai_0 _22884_ (.A1(_04964_),
    .A2(_05167_),
    .B1(_05179_),
    .Y(_00637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_348 ();
 sky130_fd_sc_hd__nand2_1 _22886_ (.A(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .B(_05167_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21ai_0 _22887_ (.A1(_02145_),
    .A2(_05167_),
    .B1(_05181_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _22888_ (.A(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .B(_05167_),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_0 _22889_ (.A1(_02297_),
    .A2(_05167_),
    .B1(_05182_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _22890_ (.A(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .B(_05167_),
    .Y(_05183_));
 sky130_fd_sc_hd__o21ai_0 _22891_ (.A1(_02414_),
    .A2(_05167_),
    .B1(_05183_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _22892_ (.A(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .B(_05167_),
    .Y(_05184_));
 sky130_fd_sc_hd__o21ai_0 _22893_ (.A1(_02535_),
    .A2(_05167_),
    .B1(_05184_),
    .Y(_00641_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_347 ();
 sky130_fd_sc_hd__nand2_1 _22895_ (.A(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .B(_05167_),
    .Y(_05186_));
 sky130_fd_sc_hd__o21ai_0 _22896_ (.A1(_02628_),
    .A2(_05167_),
    .B1(_05186_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_1 _22897_ (.A(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .B(_05167_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21ai_0 _22898_ (.A1(net3453),
    .A2(_05167_),
    .B1(_05187_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _22899_ (.A(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .B(_05167_),
    .Y(_05188_));
 sky130_fd_sc_hd__o21ai_0 _22900_ (.A1(_02837_),
    .A2(_05167_),
    .B1(_05188_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_1 _22901_ (.A(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .B(_05167_),
    .Y(_05189_));
 sky130_fd_sc_hd__o21ai_0 _22902_ (.A1(_02963_),
    .A2(_05167_),
    .B1(_05189_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _22903_ (.A(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .B(_05167_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21ai_0 _22904_ (.A1(net3447),
    .A2(_05167_),
    .B1(_05190_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_8 _22905_ (.A(net3828),
    .B(_05014_),
    .Y(_05191_));
 sky130_fd_sc_hd__nor2_4 _22906_ (.A(_05099_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__nand2_1 _22907_ (.A(net3446),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__nand2_1 _22908_ (.A(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .B(_05167_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_1 _22909_ (.A(_05193_),
    .B(_05194_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _22910_ (.A(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .B(_05167_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ai_0 _22911_ (.A1(net3425),
    .A2(_05167_),
    .B1(_05195_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _22912_ (.A(net3416),
    .B(_05192_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _22913_ (.A(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .B(_05167_),
    .Y(_05197_));
 sky130_fd_sc_hd__nand2_1 _22914_ (.A(_05196_),
    .B(_05197_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _22915_ (.A(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .B(_05167_),
    .Y(_05198_));
 sky130_fd_sc_hd__o21ai_0 _22916_ (.A1(net3433),
    .A2(_05167_),
    .B1(_05198_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2_1 _22917_ (.A(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .B(_05167_),
    .Y(_05199_));
 sky130_fd_sc_hd__o21ai_0 _22918_ (.A1(net3413),
    .A2(_05167_),
    .B1(_05199_),
    .Y(_00651_));
 sky130_fd_sc_hd__mux2_1 _22919_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A1(net3412),
    .S(_05192_),
    .X(_00652_));
 sky130_fd_sc_hd__nand2_1 _22920_ (.A(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .B(_05167_),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ai_0 _22921_ (.A1(net3411),
    .A2(_05167_),
    .B1(_05200_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _22922_ (.A(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .B(_05167_),
    .Y(_05201_));
 sky130_fd_sc_hd__o21ai_0 _22923_ (.A1(net3410),
    .A2(_05167_),
    .B1(_05201_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _22924_ (.A(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .B(_05167_),
    .Y(_05202_));
 sky130_fd_sc_hd__o21ai_0 _22925_ (.A1(net3409),
    .A2(_05167_),
    .B1(_05202_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _22926_ (.A(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .B(_05167_),
    .Y(_05203_));
 sky130_fd_sc_hd__o21ai_0 _22927_ (.A1(net3408),
    .A2(_05167_),
    .B1(_05203_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _22928_ (.A(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .B(_05167_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21ai_0 _22929_ (.A1(net3407),
    .A2(_05167_),
    .B1(_05204_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _22930_ (.A(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .B(_05167_),
    .Y(_05205_));
 sky130_fd_sc_hd__o21ai_0 _22931_ (.A1(net3406),
    .A2(_05167_),
    .B1(_05205_),
    .Y(_00658_));
 sky130_fd_sc_hd__nor2_1 _22932_ (.A(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .B(_05192_),
    .Y(_05206_));
 sky130_fd_sc_hd__a31oi_1 _22933_ (.A1(net3405),
    .A2(net3457),
    .A3(_05192_),
    .B1(_05206_),
    .Y(_00659_));
 sky130_fd_sc_hd__mux2_1 _22934_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A1(net3404),
    .S(_05192_),
    .X(_00660_));
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_04920_),
    .B(_05167_),
    .Y(_05207_));
 sky130_fd_sc_hd__a22o_1 _22936_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A2(_05167_),
    .B1(_05207_),
    .B2(net3403),
    .X(_00661_));
 sky130_fd_sc_hd__nand2_8 _22937_ (.A(_02151_),
    .B(_05013_),
    .Y(_05208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_344 ();
 sky130_fd_sc_hd__nand2_1 _22941_ (.A(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .B(_05208_),
    .Y(_05212_));
 sky130_fd_sc_hd__o21ai_0 _22942_ (.A1(_05011_),
    .A2(_05208_),
    .B1(_05212_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _22943_ (.A(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .B(_05208_),
    .Y(_05213_));
 sky130_fd_sc_hd__o21ai_0 _22944_ (.A1(_05039_),
    .A2(_05208_),
    .B1(_05213_),
    .Y(_00663_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_343 ();
 sky130_fd_sc_hd__nand2_1 _22946_ (.A(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .B(_05208_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21ai_0 _22947_ (.A1(_05059_),
    .A2(_05208_),
    .B1(_05215_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _22948_ (.A(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .B(_05208_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21ai_0 _22949_ (.A1(net3463),
    .A2(_05208_),
    .B1(_05216_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _22950_ (.A(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .B(_05208_),
    .Y(_05217_));
 sky130_fd_sc_hd__o21ai_0 _22951_ (.A1(net3459),
    .A2(_05208_),
    .B1(_05217_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _22952_ (.A(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .B(_05208_),
    .Y(_05218_));
 sky130_fd_sc_hd__o21ai_0 _22953_ (.A1(_04483_),
    .A2(_05208_),
    .B1(_05218_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _22954_ (.A(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .B(_05208_),
    .Y(_05219_));
 sky130_fd_sc_hd__o21ai_0 _22955_ (.A1(net3444),
    .A2(_05208_),
    .B1(_05219_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _22956_ (.A(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .B(_05208_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ai_0 _22957_ (.A1(_04964_),
    .A2(_05208_),
    .B1(_05220_),
    .Y(_00669_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_342 ();
 sky130_fd_sc_hd__nand2_1 _22959_ (.A(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .B(_05208_),
    .Y(_05222_));
 sky130_fd_sc_hd__o21ai_0 _22960_ (.A1(_02145_),
    .A2(_05208_),
    .B1(_05222_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _22961_ (.A(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .B(_05208_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_0 _22962_ (.A1(_02297_),
    .A2(_05208_),
    .B1(_05223_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _22963_ (.A(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .B(_05208_),
    .Y(_05224_));
 sky130_fd_sc_hd__o21ai_0 _22964_ (.A1(_02414_),
    .A2(_05208_),
    .B1(_05224_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _22965_ (.A(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .B(_05208_),
    .Y(_05225_));
 sky130_fd_sc_hd__o21ai_0 _22966_ (.A1(_02535_),
    .A2(_05208_),
    .B1(_05225_),
    .Y(_00673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_341 ();
 sky130_fd_sc_hd__nand2_1 _22968_ (.A(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .B(_05208_),
    .Y(_05227_));
 sky130_fd_sc_hd__o21ai_0 _22969_ (.A1(_02628_),
    .A2(_05208_),
    .B1(_05227_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _22970_ (.A(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .B(_05208_),
    .Y(_05228_));
 sky130_fd_sc_hd__o21ai_0 _22971_ (.A1(net3453),
    .A2(_05208_),
    .B1(_05228_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .B(_05208_),
    .Y(_05229_));
 sky130_fd_sc_hd__o21ai_0 _22973_ (.A1(_02837_),
    .A2(_05208_),
    .B1(_05229_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _22974_ (.A(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .B(_05208_),
    .Y(_05230_));
 sky130_fd_sc_hd__o21ai_0 _22975_ (.A1(_02963_),
    .A2(_05208_),
    .B1(_05230_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _22976_ (.A(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .B(_05208_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21ai_0 _22977_ (.A1(net3447),
    .A2(_05208_),
    .B1(_05231_),
    .Y(_00678_));
 sky130_fd_sc_hd__nor2_4 _22978_ (.A(_03094_),
    .B(_05099_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand2_1 _22979_ (.A(net3446),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _22980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .B(_05208_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_1 _22981_ (.A(_05233_),
    .B(_05234_),
    .Y(_00679_));
 sky130_fd_sc_hd__nand2_1 _22982_ (.A(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .B(_05208_),
    .Y(_05235_));
 sky130_fd_sc_hd__o21ai_0 _22983_ (.A1(net3425),
    .A2(_05208_),
    .B1(_05235_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _22984_ (.A(net3416),
    .B(_05232_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _22985_ (.A(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .B(_05208_),
    .Y(_05237_));
 sky130_fd_sc_hd__nand2_1 _22986_ (.A(_05236_),
    .B(_05237_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand2_1 _22987_ (.A(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .B(_05208_),
    .Y(_05238_));
 sky130_fd_sc_hd__o21ai_0 _22988_ (.A1(net3433),
    .A2(_05208_),
    .B1(_05238_),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_1 _22989_ (.A(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .B(_05208_),
    .Y(_05239_));
 sky130_fd_sc_hd__o21ai_0 _22990_ (.A1(net3413),
    .A2(_05208_),
    .B1(_05239_),
    .Y(_00683_));
 sky130_fd_sc_hd__mux2_1 _22991_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .A1(net3412),
    .S(_05232_),
    .X(_00684_));
 sky130_fd_sc_hd__nand2_1 _22992_ (.A(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .B(_05208_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ai_0 _22993_ (.A1(net3411),
    .A2(_05208_),
    .B1(_05240_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_1 _22994_ (.A(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .B(_05208_),
    .Y(_05241_));
 sky130_fd_sc_hd__o21ai_0 _22995_ (.A1(net3410),
    .A2(_05208_),
    .B1(_05241_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _22996_ (.A(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .B(_05208_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21ai_0 _22997_ (.A1(net3409),
    .A2(_05208_),
    .B1(_05242_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _22998_ (.A(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .B(_05208_),
    .Y(_05243_));
 sky130_fd_sc_hd__o21ai_0 _22999_ (.A1(net3408),
    .A2(_05208_),
    .B1(_05243_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _23000_ (.A(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .B(_05208_),
    .Y(_05244_));
 sky130_fd_sc_hd__o21ai_0 _23001_ (.A1(net3407),
    .A2(_05208_),
    .B1(_05244_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _23002_ (.A(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .B(_05208_),
    .Y(_05245_));
 sky130_fd_sc_hd__o21ai_0 _23003_ (.A1(net3406),
    .A2(_05208_),
    .B1(_05245_),
    .Y(_00690_));
 sky130_fd_sc_hd__nor2_1 _23004_ (.A(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .B(_05232_),
    .Y(_05246_));
 sky130_fd_sc_hd__a31oi_1 _23005_ (.A1(net3405),
    .A2(net3457),
    .A3(_05232_),
    .B1(_05246_),
    .Y(_00691_));
 sky130_fd_sc_hd__mux2_1 _23006_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .A1(net3404),
    .S(_05232_),
    .X(_00692_));
 sky130_fd_sc_hd__nor2_1 _23007_ (.A(_04920_),
    .B(_05208_),
    .Y(_05247_));
 sky130_fd_sc_hd__a22o_1 _23008_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .A2(_05208_),
    .B1(_05247_),
    .B2(net3403),
    .X(_00693_));
 sky130_fd_sc_hd__nor3b_4 _23009_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .C_N(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Y(_05248_));
 sky130_fd_sc_hd__nand2_8 _23010_ (.A(_05015_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_338 ();
 sky130_fd_sc_hd__nand2_1 _23014_ (.A(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .B(_05249_),
    .Y(_05253_));
 sky130_fd_sc_hd__o21ai_0 _23015_ (.A1(_05011_),
    .A2(_05249_),
    .B1(_05253_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_1 _23016_ (.A(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .B(_05249_),
    .Y(_05254_));
 sky130_fd_sc_hd__o21ai_0 _23017_ (.A1(_05039_),
    .A2(_05249_),
    .B1(_05254_),
    .Y(_00695_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_337 ();
 sky130_fd_sc_hd__nand2_1 _23019_ (.A(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .B(_05249_),
    .Y(_05256_));
 sky130_fd_sc_hd__o21ai_0 _23020_ (.A1(_05059_),
    .A2(_05249_),
    .B1(_05256_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _23021_ (.A(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .B(_05249_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21ai_0 _23022_ (.A1(net3463),
    .A2(_05249_),
    .B1(_05257_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _23023_ (.A(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .B(_05249_),
    .Y(_05258_));
 sky130_fd_sc_hd__o21ai_0 _23024_ (.A1(net3459),
    .A2(_05249_),
    .B1(_05258_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _23025_ (.A(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .B(_05249_),
    .Y(_05259_));
 sky130_fd_sc_hd__o21ai_0 _23026_ (.A1(_04483_),
    .A2(_05249_),
    .B1(_05259_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _23027_ (.A(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .B(_05249_),
    .Y(_05260_));
 sky130_fd_sc_hd__o21ai_0 _23028_ (.A1(net3444),
    .A2(_05249_),
    .B1(_05260_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _23029_ (.A(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .B(_05249_),
    .Y(_05261_));
 sky130_fd_sc_hd__o21ai_0 _23030_ (.A1(_04964_),
    .A2(_05249_),
    .B1(_05261_),
    .Y(_00701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_336 ();
 sky130_fd_sc_hd__nand2_1 _23032_ (.A(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .B(_05249_),
    .Y(_05263_));
 sky130_fd_sc_hd__o21ai_0 _23033_ (.A1(_02145_),
    .A2(_05249_),
    .B1(_05263_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _23034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .B(_05249_),
    .Y(_05264_));
 sky130_fd_sc_hd__o21ai_0 _23035_ (.A1(_02297_),
    .A2(_05249_),
    .B1(_05264_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _23036_ (.A(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .B(_05249_),
    .Y(_05265_));
 sky130_fd_sc_hd__o21ai_0 _23037_ (.A1(_02414_),
    .A2(_05249_),
    .B1(_05265_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _23038_ (.A(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .B(_05249_),
    .Y(_05266_));
 sky130_fd_sc_hd__o21ai_0 _23039_ (.A1(_02535_),
    .A2(_05249_),
    .B1(_05266_),
    .Y(_00705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_335 ();
 sky130_fd_sc_hd__nand2_1 _23041_ (.A(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .B(_05249_),
    .Y(_05268_));
 sky130_fd_sc_hd__o21ai_0 _23042_ (.A1(_02628_),
    .A2(_05249_),
    .B1(_05268_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .B(_05249_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_0 _23044_ (.A1(net3453),
    .A2(_05249_),
    .B1(_05269_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand2_1 _23045_ (.A(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .B(_05249_),
    .Y(_05270_));
 sky130_fd_sc_hd__o21ai_0 _23046_ (.A1(_02837_),
    .A2(_05249_),
    .B1(_05270_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _23047_ (.A(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .B(_05249_),
    .Y(_05271_));
 sky130_fd_sc_hd__o21ai_0 _23048_ (.A1(_02963_),
    .A2(_05249_),
    .B1(_05271_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _23049_ (.A(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .B(_05249_),
    .Y(_05272_));
 sky130_fd_sc_hd__o21ai_0 _23050_ (.A1(net3447),
    .A2(_05249_),
    .B1(_05272_),
    .Y(_00710_));
 sky130_fd_sc_hd__or3b_4 _23051_ (.A(net3827),
    .B(net3945),
    .C_N(net3946),
    .X(_05273_));
 sky130_fd_sc_hd__nor2_4 _23052_ (.A(_05100_),
    .B(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _23053_ (.A(net3446),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _23054_ (.A(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .B(_05249_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_1 _23055_ (.A(_05275_),
    .B(_05276_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _23056_ (.A(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .B(_05249_),
    .Y(_05277_));
 sky130_fd_sc_hd__o21ai_0 _23057_ (.A1(net3425),
    .A2(_05249_),
    .B1(_05277_),
    .Y(_00712_));
 sky130_fd_sc_hd__nand2_1 _23058_ (.A(net3416),
    .B(_05274_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_1 _23059_ (.A(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .B(_05249_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _23060_ (.A(_05278_),
    .B(_05279_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _23061_ (.A(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .B(_05249_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21ai_0 _23062_ (.A1(net3433),
    .A2(_05249_),
    .B1(_05280_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _23063_ (.A(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .B(_05249_),
    .Y(_05281_));
 sky130_fd_sc_hd__o21ai_0 _23064_ (.A1(net3413),
    .A2(_05249_),
    .B1(_05281_),
    .Y(_00715_));
 sky130_fd_sc_hd__mux2_1 _23065_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(net3412),
    .S(_05274_),
    .X(_00716_));
 sky130_fd_sc_hd__nand2_1 _23066_ (.A(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .B(_05249_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21ai_0 _23067_ (.A1(net3411),
    .A2(_05249_),
    .B1(_05282_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand2_1 _23068_ (.A(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .B(_05249_),
    .Y(_05283_));
 sky130_fd_sc_hd__o21ai_0 _23069_ (.A1(net3410),
    .A2(_05249_),
    .B1(_05283_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _23070_ (.A(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .B(_05249_),
    .Y(_05284_));
 sky130_fd_sc_hd__o21ai_0 _23071_ (.A1(net3409),
    .A2(_05249_),
    .B1(_05284_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_1 _23072_ (.A(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .B(_05249_),
    .Y(_05285_));
 sky130_fd_sc_hd__o21ai_0 _23073_ (.A1(net3408),
    .A2(_05249_),
    .B1(_05285_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_1 _23074_ (.A(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .B(_05249_),
    .Y(_05286_));
 sky130_fd_sc_hd__o21ai_0 _23075_ (.A1(net3407),
    .A2(_05249_),
    .B1(_05286_),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_1 _23076_ (.A(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .B(_05249_),
    .Y(_05287_));
 sky130_fd_sc_hd__o21ai_0 _23077_ (.A1(net3406),
    .A2(_05249_),
    .B1(_05287_),
    .Y(_00722_));
 sky130_fd_sc_hd__nor2_1 _23078_ (.A(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .B(_05274_),
    .Y(_05288_));
 sky130_fd_sc_hd__a31oi_1 _23079_ (.A1(net3405),
    .A2(net3457),
    .A3(_05274_),
    .B1(_05288_),
    .Y(_00723_));
 sky130_fd_sc_hd__mux2_1 _23080_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(net3404),
    .S(_05274_),
    .X(_00724_));
 sky130_fd_sc_hd__nor2_1 _23081_ (.A(_04920_),
    .B(_05249_),
    .Y(_05289_));
 sky130_fd_sc_hd__a22o_1 _23082_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A2(_05249_),
    .B1(_05289_),
    .B2(net3403),
    .X(_00725_));
 sky130_fd_sc_hd__nand2_8 _23083_ (.A(_05122_),
    .B(_05248_),
    .Y(_05290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_332 ();
 sky130_fd_sc_hd__nand2_1 _23087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .B(_05290_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21ai_0 _23088_ (.A1(_05011_),
    .A2(_05290_),
    .B1(_05294_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_1 _23089_ (.A(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .B(_05290_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_0 _23090_ (.A1(_05039_),
    .A2(_05290_),
    .B1(_05295_),
    .Y(_00727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_331 ();
 sky130_fd_sc_hd__nand2_1 _23092_ (.A(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .B(_05290_),
    .Y(_05297_));
 sky130_fd_sc_hd__o21ai_0 _23093_ (.A1(_05059_),
    .A2(_05290_),
    .B1(_05297_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _23094_ (.A(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .B(_05290_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ai_0 _23095_ (.A1(net3463),
    .A2(_05290_),
    .B1(_05298_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _23096_ (.A(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .B(_05290_),
    .Y(_05299_));
 sky130_fd_sc_hd__o21ai_0 _23097_ (.A1(net3459),
    .A2(_05290_),
    .B1(_05299_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _23098_ (.A(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .B(_05290_),
    .Y(_05300_));
 sky130_fd_sc_hd__o21ai_0 _23099_ (.A1(_04483_),
    .A2(_05290_),
    .B1(_05300_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _23100_ (.A(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .B(_05290_),
    .Y(_05301_));
 sky130_fd_sc_hd__o21ai_0 _23101_ (.A1(net3444),
    .A2(_05290_),
    .B1(_05301_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _23102_ (.A(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .B(_05290_),
    .Y(_05302_));
 sky130_fd_sc_hd__o21ai_0 _23103_ (.A1(_04964_),
    .A2(_05290_),
    .B1(_05302_),
    .Y(_00733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_330 ();
 sky130_fd_sc_hd__nand2_1 _23105_ (.A(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .B(_05290_),
    .Y(_05304_));
 sky130_fd_sc_hd__o21ai_0 _23106_ (.A1(_02145_),
    .A2(_05290_),
    .B1(_05304_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _23107_ (.A(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .B(_05290_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21ai_0 _23108_ (.A1(_02297_),
    .A2(_05290_),
    .B1(_05305_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand2_1 _23109_ (.A(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .B(_05290_),
    .Y(_05306_));
 sky130_fd_sc_hd__o21ai_0 _23110_ (.A1(_02414_),
    .A2(_05290_),
    .B1(_05306_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _23111_ (.A(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .B(_05290_),
    .Y(_05307_));
 sky130_fd_sc_hd__o21ai_0 _23112_ (.A1(_02535_),
    .A2(_05290_),
    .B1(_05307_),
    .Y(_00737_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_329 ();
 sky130_fd_sc_hd__nand2_1 _23114_ (.A(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .B(_05290_),
    .Y(_05309_));
 sky130_fd_sc_hd__o21ai_0 _23115_ (.A1(_02628_),
    .A2(_05290_),
    .B1(_05309_),
    .Y(_00738_));
 sky130_fd_sc_hd__nand2_1 _23116_ (.A(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .B(_05290_),
    .Y(_05310_));
 sky130_fd_sc_hd__o21ai_0 _23117_ (.A1(net3453),
    .A2(_05290_),
    .B1(_05310_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _23118_ (.A(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .B(_05290_),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_0 _23119_ (.A1(_02837_),
    .A2(_05290_),
    .B1(_05311_),
    .Y(_00740_));
 sky130_fd_sc_hd__nand2_1 _23120_ (.A(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .B(_05290_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_0 _23121_ (.A1(_02963_),
    .A2(_05290_),
    .B1(_05312_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand2_1 _23122_ (.A(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .B(_05290_),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_0 _23123_ (.A1(net3447),
    .A2(_05290_),
    .B1(_05313_),
    .Y(_00742_));
 sky130_fd_sc_hd__nor2_4 _23124_ (.A(_05147_),
    .B(_05273_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand2_1 _23125_ (.A(net3446),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .B(_05290_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _23127_ (.A(_05315_),
    .B(_05316_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _23128_ (.A(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .B(_05290_),
    .Y(_05317_));
 sky130_fd_sc_hd__o21ai_0 _23129_ (.A1(net3425),
    .A2(_05290_),
    .B1(_05317_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_1 _23130_ (.A(net3416),
    .B(_05314_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _23131_ (.A(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .B(_05290_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_1 _23132_ (.A(_05318_),
    .B(_05319_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _23133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .B(_05290_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21ai_0 _23134_ (.A1(net3433),
    .A2(_05290_),
    .B1(_05320_),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _23135_ (.A(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .B(_05290_),
    .Y(_05321_));
 sky130_fd_sc_hd__o21ai_0 _23136_ (.A1(net3413),
    .A2(_05290_),
    .B1(_05321_),
    .Y(_00747_));
 sky130_fd_sc_hd__mux2_1 _23137_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A1(net3412),
    .S(_05314_),
    .X(_00748_));
 sky130_fd_sc_hd__nand2_1 _23138_ (.A(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .B(_05290_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_0 _23139_ (.A1(net3411),
    .A2(_05290_),
    .B1(_05322_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _23140_ (.A(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .B(_05290_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21ai_0 _23141_ (.A1(net3410),
    .A2(_05290_),
    .B1(_05323_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand2_1 _23142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .B(_05290_),
    .Y(_05324_));
 sky130_fd_sc_hd__o21ai_0 _23143_ (.A1(net3409),
    .A2(_05290_),
    .B1(_05324_),
    .Y(_00751_));
 sky130_fd_sc_hd__nand2_1 _23144_ (.A(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .B(_05290_),
    .Y(_05325_));
 sky130_fd_sc_hd__o21ai_0 _23145_ (.A1(net3408),
    .A2(_05290_),
    .B1(_05325_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand2_1 _23146_ (.A(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .B(_05290_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_0 _23147_ (.A1(net3407),
    .A2(_05290_),
    .B1(_05326_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _23148_ (.A(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .B(_05290_),
    .Y(_05327_));
 sky130_fd_sc_hd__o21ai_0 _23149_ (.A1(net3406),
    .A2(_05290_),
    .B1(_05327_),
    .Y(_00754_));
 sky130_fd_sc_hd__nor2_1 _23150_ (.A(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .B(_05314_),
    .Y(_05328_));
 sky130_fd_sc_hd__a31oi_1 _23151_ (.A1(net3405),
    .A2(net3457),
    .A3(_05314_),
    .B1(_05328_),
    .Y(_00755_));
 sky130_fd_sc_hd__mux2_1 _23152_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A1(net3404),
    .S(_05314_),
    .X(_00756_));
 sky130_fd_sc_hd__nor2_1 _23153_ (.A(_04920_),
    .B(_05290_),
    .Y(_05329_));
 sky130_fd_sc_hd__a22o_1 _23154_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A2(_05290_),
    .B1(_05329_),
    .B2(net3403),
    .X(_00757_));
 sky130_fd_sc_hd__nand2_8 _23155_ (.A(_05165_),
    .B(_05248_),
    .Y(_05330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_326 ();
 sky130_fd_sc_hd__nand2_1 _23159_ (.A(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .B(_05330_),
    .Y(_05334_));
 sky130_fd_sc_hd__o21ai_0 _23160_ (.A1(_05011_),
    .A2(_05330_),
    .B1(_05334_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand2_1 _23161_ (.A(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .B(_05330_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21ai_0 _23162_ (.A1(_05039_),
    .A2(_05330_),
    .B1(_05335_),
    .Y(_00759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_325 ();
 sky130_fd_sc_hd__nand2_1 _23164_ (.A(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .B(_05330_),
    .Y(_05337_));
 sky130_fd_sc_hd__o21ai_0 _23165_ (.A1(_05059_),
    .A2(_05330_),
    .B1(_05337_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand2_1 _23166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .B(_05330_),
    .Y(_05338_));
 sky130_fd_sc_hd__o21ai_0 _23167_ (.A1(net3463),
    .A2(_05330_),
    .B1(_05338_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _23168_ (.A(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .B(_05330_),
    .Y(_05339_));
 sky130_fd_sc_hd__o21ai_0 _23169_ (.A1(net3459),
    .A2(_05330_),
    .B1(_05339_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _23170_ (.A(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .B(_05330_),
    .Y(_05340_));
 sky130_fd_sc_hd__o21ai_0 _23171_ (.A1(_04483_),
    .A2(_05330_),
    .B1(_05340_),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _23172_ (.A(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .B(_05330_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21ai_0 _23173_ (.A1(net3444),
    .A2(_05330_),
    .B1(_05341_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _23174_ (.A(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .B(_05330_),
    .Y(_05342_));
 sky130_fd_sc_hd__o21ai_0 _23175_ (.A1(_04964_),
    .A2(_05330_),
    .B1(_05342_),
    .Y(_00765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_324 ();
 sky130_fd_sc_hd__nand2_1 _23177_ (.A(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .B(_05330_),
    .Y(_05344_));
 sky130_fd_sc_hd__o21ai_0 _23178_ (.A1(_02145_),
    .A2(_05330_),
    .B1(_05344_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _23179_ (.A(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .B(_05330_),
    .Y(_05345_));
 sky130_fd_sc_hd__o21ai_0 _23180_ (.A1(_02297_),
    .A2(_05330_),
    .B1(_05345_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_8 _23181_ (.A(_10519_),
    .B(net3455),
    .Y(_05346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_321 ();
 sky130_fd_sc_hd__nand2_1 _23185_ (.A(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B(_05346_),
    .Y(_05350_));
 sky130_fd_sc_hd__o21ai_0 _23186_ (.A1(_05011_),
    .A2(_05346_),
    .B1(_05350_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _23187_ (.A(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .B(_05330_),
    .Y(_05351_));
 sky130_fd_sc_hd__o21ai_0 _23188_ (.A1(_02414_),
    .A2(_05330_),
    .B1(_05351_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _23189_ (.A(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .B(_05330_),
    .Y(_05352_));
 sky130_fd_sc_hd__o21ai_0 _23190_ (.A1(_02535_),
    .A2(_05330_),
    .B1(_05352_),
    .Y(_00770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_320 ();
 sky130_fd_sc_hd__nand2_1 _23192_ (.A(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .B(_05330_),
    .Y(_05354_));
 sky130_fd_sc_hd__o21ai_0 _23193_ (.A1(_02628_),
    .A2(_05330_),
    .B1(_05354_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _23194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .B(_05330_),
    .Y(_05355_));
 sky130_fd_sc_hd__o21ai_0 _23195_ (.A1(net3453),
    .A2(_05330_),
    .B1(_05355_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand2_1 _23196_ (.A(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .B(_05330_),
    .Y(_05356_));
 sky130_fd_sc_hd__o21ai_0 _23197_ (.A1(_02837_),
    .A2(_05330_),
    .B1(_05356_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_1 _23198_ (.A(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .B(_05330_),
    .Y(_05357_));
 sky130_fd_sc_hd__o21ai_0 _23199_ (.A1(_02963_),
    .A2(_05330_),
    .B1(_05357_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _23200_ (.A(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .B(_05330_),
    .Y(_05358_));
 sky130_fd_sc_hd__o21ai_0 _23201_ (.A1(net3447),
    .A2(_05330_),
    .B1(_05358_),
    .Y(_00775_));
 sky130_fd_sc_hd__nor2_4 _23202_ (.A(_05191_),
    .B(_05273_),
    .Y(_05359_));
 sky130_fd_sc_hd__nand2_1 _23203_ (.A(net3446),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _23204_ (.A(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .B(_05330_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _23205_ (.A(_05360_),
    .B(_05361_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _23206_ (.A(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .B(_05330_),
    .Y(_05362_));
 sky130_fd_sc_hd__o21ai_0 _23207_ (.A1(net3425),
    .A2(_05330_),
    .B1(_05362_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _23208_ (.A(net3416),
    .B(_05359_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _23209_ (.A(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .B(_05330_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _23210_ (.A(_05363_),
    .B(_05364_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _23211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .B(_05346_),
    .Y(_05365_));
 sky130_fd_sc_hd__o21ai_0 _23212_ (.A1(_05039_),
    .A2(_05346_),
    .B1(_05365_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_1 _23213_ (.A(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .B(_05330_),
    .Y(_05366_));
 sky130_fd_sc_hd__o21ai_0 _23214_ (.A1(net3433),
    .A2(_05330_),
    .B1(_05366_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _23215_ (.A(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .B(_05330_),
    .Y(_05367_));
 sky130_fd_sc_hd__o21ai_0 _23216_ (.A1(net3413),
    .A2(_05330_),
    .B1(_05367_),
    .Y(_00781_));
 sky130_fd_sc_hd__mux2_1 _23217_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A1(net3412),
    .S(_05359_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .B(_05330_),
    .Y(_05368_));
 sky130_fd_sc_hd__o21ai_0 _23219_ (.A1(net3411),
    .A2(_05330_),
    .B1(_05368_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand2_1 _23220_ (.A(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .B(_05330_),
    .Y(_05369_));
 sky130_fd_sc_hd__o21ai_0 _23221_ (.A1(net3410),
    .A2(_05330_),
    .B1(_05369_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _23222_ (.A(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .B(_05330_),
    .Y(_05370_));
 sky130_fd_sc_hd__o21ai_0 _23223_ (.A1(net3409),
    .A2(_05330_),
    .B1(_05370_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand2_1 _23224_ (.A(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .B(_05330_),
    .Y(_05371_));
 sky130_fd_sc_hd__o21ai_0 _23225_ (.A1(net3408),
    .A2(_05330_),
    .B1(_05371_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_1 _23226_ (.A(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .B(_05330_),
    .Y(_05372_));
 sky130_fd_sc_hd__o21ai_0 _23227_ (.A1(net3407),
    .A2(_05330_),
    .B1(_05372_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_1 _23228_ (.A(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .B(_05330_),
    .Y(_05373_));
 sky130_fd_sc_hd__o21ai_0 _23229_ (.A1(net3406),
    .A2(_05330_),
    .B1(_05373_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor2_1 _23230_ (.A(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .B(_05359_),
    .Y(_05374_));
 sky130_fd_sc_hd__a31oi_1 _23231_ (.A1(net3405),
    .A2(net3457),
    .A3(_05359_),
    .B1(_05374_),
    .Y(_00789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_319 ();
 sky130_fd_sc_hd__nand2_1 _23233_ (.A(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .B(_05346_),
    .Y(_05376_));
 sky130_fd_sc_hd__o21ai_0 _23234_ (.A1(_05059_),
    .A2(_05346_),
    .B1(_05376_),
    .Y(_00790_));
 sky130_fd_sc_hd__mux2_1 _23235_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A1(net3404),
    .S(_05359_),
    .X(_00791_));
 sky130_fd_sc_hd__nor2_1 _23236_ (.A(net3464),
    .B(_05330_),
    .Y(_05377_));
 sky130_fd_sc_hd__a22o_1 _23237_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A2(_05330_),
    .B1(_05377_),
    .B2(net3403),
    .X(_00792_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_318 ();
 sky130_fd_sc_hd__nand2_8 _23239_ (.A(_02151_),
    .B(_05248_),
    .Y(_05379_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_315 ();
 sky130_fd_sc_hd__nand2_1 _23243_ (.A(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .B(_05379_),
    .Y(_05383_));
 sky130_fd_sc_hd__o21ai_0 _23244_ (.A1(_05011_),
    .A2(_05379_),
    .B1(_05383_),
    .Y(_00793_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_314 ();
 sky130_fd_sc_hd__nand2_1 _23246_ (.A(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .B(_05379_),
    .Y(_05385_));
 sky130_fd_sc_hd__o21ai_0 _23247_ (.A1(_05039_),
    .A2(_05379_),
    .B1(_05385_),
    .Y(_00794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_312 ();
 sky130_fd_sc_hd__nand2_1 _23250_ (.A(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .B(_05379_),
    .Y(_05388_));
 sky130_fd_sc_hd__o21ai_0 _23251_ (.A1(_05059_),
    .A2(_05379_),
    .B1(_05388_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _23252_ (.A(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .B(_05379_),
    .Y(_05389_));
 sky130_fd_sc_hd__o21ai_0 _23253_ (.A1(net3463),
    .A2(_05379_),
    .B1(_05389_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand2_1 _23254_ (.A(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .B(_05379_),
    .Y(_05390_));
 sky130_fd_sc_hd__o21ai_0 _23255_ (.A1(net3459),
    .A2(_05379_),
    .B1(_05390_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _23256_ (.A(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .B(_05379_),
    .Y(_05391_));
 sky130_fd_sc_hd__o21ai_0 _23257_ (.A1(_04483_),
    .A2(_05379_),
    .B1(_05391_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _23258_ (.A(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .B(_05379_),
    .Y(_05392_));
 sky130_fd_sc_hd__o21ai_0 _23259_ (.A1(net3444),
    .A2(_05379_),
    .B1(_05392_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _23260_ (.A(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .B(_05379_),
    .Y(_05393_));
 sky130_fd_sc_hd__o21ai_0 _23261_ (.A1(_04964_),
    .A2(_05379_),
    .B1(_05393_),
    .Y(_00800_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_311 ();
 sky130_fd_sc_hd__nand2_1 _23263_ (.A(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .B(_05346_),
    .Y(_05395_));
 sky130_fd_sc_hd__o21ai_0 _23264_ (.A1(net3463),
    .A2(_05346_),
    .B1(_05395_),
    .Y(_00801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_310 ();
 sky130_fd_sc_hd__nand2_1 _23266_ (.A(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .B(_05379_),
    .Y(_05397_));
 sky130_fd_sc_hd__o21ai_0 _23267_ (.A1(_02145_),
    .A2(_05379_),
    .B1(_05397_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand2_1 _23268_ (.A(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .B(_05379_),
    .Y(_05398_));
 sky130_fd_sc_hd__o21ai_0 _23269_ (.A1(_02297_),
    .A2(_05379_),
    .B1(_05398_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_1 _23270_ (.A(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .B(_05379_),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_0 _23271_ (.A1(_02414_),
    .A2(_05379_),
    .B1(_05399_),
    .Y(_00804_));
 sky130_fd_sc_hd__nand2_1 _23272_ (.A(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .B(_05379_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_0 _23273_ (.A1(_02535_),
    .A2(_05379_),
    .B1(_05400_),
    .Y(_00805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_309 ();
 sky130_fd_sc_hd__nand2_1 _23275_ (.A(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .B(_05379_),
    .Y(_05402_));
 sky130_fd_sc_hd__o21ai_0 _23276_ (.A1(_02628_),
    .A2(_05379_),
    .B1(_05402_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _23277_ (.A(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .B(_05379_),
    .Y(_05403_));
 sky130_fd_sc_hd__o21ai_0 _23278_ (.A1(net3453),
    .A2(_05379_),
    .B1(_05403_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_1 _23279_ (.A(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .B(_05379_),
    .Y(_05404_));
 sky130_fd_sc_hd__o21ai_0 _23280_ (.A1(_02837_),
    .A2(_05379_),
    .B1(_05404_),
    .Y(_00808_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .B(_05379_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ai_0 _23282_ (.A1(_02963_),
    .A2(_05379_),
    .B1(_05405_),
    .Y(_00809_));
 sky130_fd_sc_hd__nand2_1 _23283_ (.A(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .B(_05379_),
    .Y(_05406_));
 sky130_fd_sc_hd__o21ai_0 _23284_ (.A1(net3447),
    .A2(_05379_),
    .B1(_05406_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor2_4 _23285_ (.A(_03094_),
    .B(_05273_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _23286_ (.A(net3446),
    .B(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _23287_ (.A(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .B(_05379_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _23288_ (.A(_05408_),
    .B(_05409_),
    .Y(_00811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_308 ();
 sky130_fd_sc_hd__nand2_1 _23290_ (.A(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B(_05346_),
    .Y(_05411_));
 sky130_fd_sc_hd__o21ai_0 _23291_ (.A1(net3459),
    .A2(_05346_),
    .B1(_05411_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _23292_ (.A(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .B(_05379_),
    .Y(_05412_));
 sky130_fd_sc_hd__o21ai_0 _23293_ (.A1(net3425),
    .A2(_05379_),
    .B1(_05412_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _23294_ (.A(net3416),
    .B(_05407_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _23295_ (.A(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .B(_05379_),
    .Y(_05414_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_05413_),
    .B(_05414_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _23297_ (.A(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .B(_05379_),
    .Y(_05415_));
 sky130_fd_sc_hd__o21ai_0 _23298_ (.A1(net3433),
    .A2(_05379_),
    .B1(_05415_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _23299_ (.A(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .B(_05379_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21ai_0 _23300_ (.A1(net3413),
    .A2(_05379_),
    .B1(_05416_),
    .Y(_00816_));
 sky130_fd_sc_hd__mux2_1 _23301_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .A1(net3412),
    .S(_05407_),
    .X(_00817_));
 sky130_fd_sc_hd__nand2_1 _23302_ (.A(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .B(_05379_),
    .Y(_05417_));
 sky130_fd_sc_hd__o21ai_0 _23303_ (.A1(net3411),
    .A2(_05379_),
    .B1(_05417_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _23304_ (.A(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .B(_05379_),
    .Y(_05418_));
 sky130_fd_sc_hd__o21ai_0 _23305_ (.A1(net3410),
    .A2(_05379_),
    .B1(_05418_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _23306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .B(_05379_),
    .Y(_05419_));
 sky130_fd_sc_hd__o21ai_0 _23307_ (.A1(net3409),
    .A2(_05379_),
    .B1(_05419_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_1 _23308_ (.A(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .B(_05379_),
    .Y(_05420_));
 sky130_fd_sc_hd__o21ai_0 _23309_ (.A1(net3408),
    .A2(_05379_),
    .B1(_05420_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _23310_ (.A(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .B(_05379_),
    .Y(_05421_));
 sky130_fd_sc_hd__o21ai_0 _23311_ (.A1(net3407),
    .A2(_05379_),
    .B1(_05421_),
    .Y(_00822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_307 ();
 sky130_fd_sc_hd__nand2_1 _23313_ (.A(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .B(_05346_),
    .Y(_05423_));
 sky130_fd_sc_hd__o21ai_0 _23314_ (.A1(_04483_),
    .A2(_05346_),
    .B1(_05423_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _23315_ (.A(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .B(_05379_),
    .Y(_05424_));
 sky130_fd_sc_hd__o21ai_0 _23316_ (.A1(net3406),
    .A2(_05379_),
    .B1(_05424_),
    .Y(_00824_));
 sky130_fd_sc_hd__nor2_1 _23317_ (.A(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .B(_05407_),
    .Y(_05425_));
 sky130_fd_sc_hd__a31oi_1 _23318_ (.A1(net3405),
    .A2(net3457),
    .A3(_05407_),
    .B1(_05425_),
    .Y(_00825_));
 sky130_fd_sc_hd__mux2_1 _23319_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .A1(net3404),
    .S(_05407_),
    .X(_00826_));
 sky130_fd_sc_hd__nor2_1 _23320_ (.A(net3464),
    .B(_05379_),
    .Y(_05426_));
 sky130_fd_sc_hd__a22o_1 _23321_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .A2(_05379_),
    .B1(_05426_),
    .B2(net3403),
    .X(_00827_));
 sky130_fd_sc_hd__nand2_2 _23322_ (.A(net3946),
    .B(net3827),
    .Y(_05427_));
 sky130_fd_sc_hd__nor2_4 _23323_ (.A(net3945),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_8 _23324_ (.A(_05015_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_304 ();
 sky130_fd_sc_hd__nand2_1 _23328_ (.A(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .B(_05429_),
    .Y(_05433_));
 sky130_fd_sc_hd__o21ai_0 _23329_ (.A1(_05011_),
    .A2(_05429_),
    .B1(_05433_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _23330_ (.A(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .B(_05429_),
    .Y(_05434_));
 sky130_fd_sc_hd__o21ai_0 _23331_ (.A1(net3456),
    .A2(_05429_),
    .B1(_05434_),
    .Y(_00829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_303 ();
 sky130_fd_sc_hd__nand2_1 _23333_ (.A(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .B(_05429_),
    .Y(_05436_));
 sky130_fd_sc_hd__o21ai_0 _23334_ (.A1(_05059_),
    .A2(_05429_),
    .B1(_05436_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _23335_ (.A(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .B(_05429_),
    .Y(_05437_));
 sky130_fd_sc_hd__o21ai_0 _23336_ (.A1(net3463),
    .A2(_05429_),
    .B1(_05437_),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .B(_05429_),
    .Y(_05438_));
 sky130_fd_sc_hd__o21ai_0 _23338_ (.A1(net3459),
    .A2(_05429_),
    .B1(_05438_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_1 _23339_ (.A(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .B(_05429_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_0 _23340_ (.A1(_04483_),
    .A2(_05429_),
    .B1(_05439_),
    .Y(_00833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_302 ();
 sky130_fd_sc_hd__nand2_1 _23342_ (.A(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .B(_05346_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21ai_0 _23343_ (.A1(net3444),
    .A2(_05346_),
    .B1(_05441_),
    .Y(_00834_));
 sky130_fd_sc_hd__nand2_1 _23344_ (.A(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .B(_05429_),
    .Y(_05442_));
 sky130_fd_sc_hd__o21ai_0 _23345_ (.A1(net3444),
    .A2(_05429_),
    .B1(_05442_),
    .Y(_00835_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_301 ();
 sky130_fd_sc_hd__nand2_1 _23347_ (.A(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .B(_05429_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_0 _23348_ (.A1(_04964_),
    .A2(_05429_),
    .B1(_05444_),
    .Y(_00836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_299 ();
 sky130_fd_sc_hd__nand2_1 _23351_ (.A(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .B(_05429_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21ai_0 _23352_ (.A1(_02145_),
    .A2(_05429_),
    .B1(_05447_),
    .Y(_00837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_298 ();
 sky130_fd_sc_hd__nand2_1 _23354_ (.A(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .B(_05429_),
    .Y(_05449_));
 sky130_fd_sc_hd__o21ai_0 _23355_ (.A1(_02297_),
    .A2(_05429_),
    .B1(_05449_),
    .Y(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_297 ();
 sky130_fd_sc_hd__nand2_1 _23357_ (.A(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .B(_05429_),
    .Y(_05451_));
 sky130_fd_sc_hd__o21ai_0 _23358_ (.A1(_02414_),
    .A2(_05429_),
    .B1(_05451_),
    .Y(_00839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_296 ();
 sky130_fd_sc_hd__nand2_1 _23360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .B(_05429_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_0 _23361_ (.A1(_02535_),
    .A2(_05429_),
    .B1(_05453_),
    .Y(_00840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_294 ();
 sky130_fd_sc_hd__nand2_1 _23364_ (.A(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .B(_05429_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_0 _23365_ (.A1(_02628_),
    .A2(_05429_),
    .B1(_05456_),
    .Y(_00841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_293 ();
 sky130_fd_sc_hd__nand2_1 _23367_ (.A(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .B(_05429_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21ai_0 _23368_ (.A1(net3453),
    .A2(_05429_),
    .B1(_05458_),
    .Y(_00842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_292 ();
 sky130_fd_sc_hd__nand2_1 _23370_ (.A(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .B(_05429_),
    .Y(_05460_));
 sky130_fd_sc_hd__o21ai_0 _23371_ (.A1(_02837_),
    .A2(_05429_),
    .B1(_05460_),
    .Y(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_291 ();
 sky130_fd_sc_hd__nand2_1 _23373_ (.A(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .B(_05429_),
    .Y(_05462_));
 sky130_fd_sc_hd__o21ai_0 _23374_ (.A1(_02963_),
    .A2(_05429_),
    .B1(_05462_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _23375_ (.A(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .B(_05346_),
    .Y(_05463_));
 sky130_fd_sc_hd__o21ai_0 _23376_ (.A1(_04964_),
    .A2(_05346_),
    .B1(_05463_),
    .Y(_00845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_290 ();
 sky130_fd_sc_hd__nand2_1 _23378_ (.A(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .B(_05429_),
    .Y(_05465_));
 sky130_fd_sc_hd__o21ai_0 _23379_ (.A1(net3447),
    .A2(_05429_),
    .B1(_05465_),
    .Y(_00846_));
 sky130_fd_sc_hd__or2_4 _23380_ (.A(net3945),
    .B(_05427_),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_4 _23381_ (.A(_05100_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _23382_ (.A(net3446),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand2_1 _23383_ (.A(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .B(_05429_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _23384_ (.A(_05468_),
    .B(_05469_),
    .Y(_00847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_289 ();
 sky130_fd_sc_hd__nand2_1 _23386_ (.A(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .B(_05429_),
    .Y(_05471_));
 sky130_fd_sc_hd__o21ai_0 _23387_ (.A1(net3425),
    .A2(_05429_),
    .B1(_05471_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand2_1 _23388_ (.A(net3416),
    .B(_05467_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _23389_ (.A(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .B(_05429_),
    .Y(_05473_));
 sky130_fd_sc_hd__nand2_1 _23390_ (.A(_05472_),
    .B(_05473_),
    .Y(_00849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_288 ();
 sky130_fd_sc_hd__nand2_1 _23392_ (.A(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .B(_05429_),
    .Y(_05475_));
 sky130_fd_sc_hd__o21ai_0 _23393_ (.A1(net3433),
    .A2(_05429_),
    .B1(_05475_),
    .Y(_00850_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_287 ();
 sky130_fd_sc_hd__nand2_1 _23395_ (.A(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .B(_05429_),
    .Y(_05477_));
 sky130_fd_sc_hd__o21ai_0 _23396_ (.A1(net3413),
    .A2(_05429_),
    .B1(_05477_),
    .Y(_00851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_286 ();
 sky130_fd_sc_hd__mux2_1 _23398_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A1(net3412),
    .S(_05467_),
    .X(_00852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_285 ();
 sky130_fd_sc_hd__nand2_1 _23400_ (.A(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .B(_05429_),
    .Y(_05480_));
 sky130_fd_sc_hd__o21ai_0 _23401_ (.A1(net3411),
    .A2(_05429_),
    .B1(_05480_),
    .Y(_00853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_284 ();
 sky130_fd_sc_hd__nand2_1 _23403_ (.A(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .B(_05429_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_0 _23404_ (.A1(net3410),
    .A2(_05429_),
    .B1(_05482_),
    .Y(_00854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_283 ();
 sky130_fd_sc_hd__nand2_1 _23406_ (.A(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .B(_05429_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_0 _23407_ (.A1(net3409),
    .A2(_05429_),
    .B1(_05484_),
    .Y(_00855_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_282 ();
 sky130_fd_sc_hd__nand2_1 _23409_ (.A(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .B(_05346_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_0 _23410_ (.A1(_02145_),
    .A2(_05346_),
    .B1(_05486_),
    .Y(_00856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_281 ();
 sky130_fd_sc_hd__nand2_1 _23412_ (.A(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .B(_05429_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21ai_0 _23413_ (.A1(net3408),
    .A2(_05429_),
    .B1(_05488_),
    .Y(_00857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_280 ();
 sky130_fd_sc_hd__nand2_1 _23415_ (.A(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .B(_05429_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_0 _23416_ (.A1(net3407),
    .A2(_05429_),
    .B1(_05490_),
    .Y(_00858_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_279 ();
 sky130_fd_sc_hd__nand2_1 _23418_ (.A(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .B(_05429_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21ai_0 _23419_ (.A1(net3406),
    .A2(_05429_),
    .B1(_05492_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor2_1 _23420_ (.A(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .B(_05467_),
    .Y(_05493_));
 sky130_fd_sc_hd__a31oi_1 _23421_ (.A1(net3405),
    .A2(net3457),
    .A3(_05467_),
    .B1(_05493_),
    .Y(_00860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_278 ();
 sky130_fd_sc_hd__mux2_1 _23423_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A1(net3404),
    .S(_05467_),
    .X(_00861_));
 sky130_fd_sc_hd__nor2_1 _23424_ (.A(_04920_),
    .B(_05429_),
    .Y(_05495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_277 ();
 sky130_fd_sc_hd__a22o_1 _23426_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A2(_05429_),
    .B1(_05495_),
    .B2(net3403),
    .X(_00862_));
 sky130_fd_sc_hd__nand2_8 _23427_ (.A(_05122_),
    .B(_05428_),
    .Y(_05497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_274 ();
 sky130_fd_sc_hd__nand2_1 _23431_ (.A(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .B(_05497_),
    .Y(_05501_));
 sky130_fd_sc_hd__o21ai_0 _23432_ (.A1(_05011_),
    .A2(_05497_),
    .B1(_05501_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand2_1 _23433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .B(_05497_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21ai_0 _23434_ (.A1(net3456),
    .A2(_05497_),
    .B1(_05502_),
    .Y(_00864_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_273 ();
 sky130_fd_sc_hd__nand2_1 _23436_ (.A(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .B(_05497_),
    .Y(_05504_));
 sky130_fd_sc_hd__o21ai_0 _23437_ (.A1(_05059_),
    .A2(_05497_),
    .B1(_05504_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _23438_ (.A(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .B(_05497_),
    .Y(_05505_));
 sky130_fd_sc_hd__o21ai_0 _23439_ (.A1(net3463),
    .A2(_05497_),
    .B1(_05505_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand2_1 _23440_ (.A(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .B(_05346_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_0 _23441_ (.A1(_02297_),
    .A2(_05346_),
    .B1(_05506_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _23442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .B(_05497_),
    .Y(_05507_));
 sky130_fd_sc_hd__o21ai_0 _23443_ (.A1(net3459),
    .A2(_05497_),
    .B1(_05507_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _23444_ (.A(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .B(_05497_),
    .Y(_05508_));
 sky130_fd_sc_hd__o21ai_0 _23445_ (.A1(_04483_),
    .A2(_05497_),
    .B1(_05508_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2_1 _23446_ (.A(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .B(_05497_),
    .Y(_05509_));
 sky130_fd_sc_hd__o21ai_0 _23447_ (.A1(net3444),
    .A2(_05497_),
    .B1(_05509_),
    .Y(_00870_));
 sky130_fd_sc_hd__nand2_1 _23448_ (.A(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .B(_05497_),
    .Y(_05510_));
 sky130_fd_sc_hd__o21ai_0 _23449_ (.A1(_04964_),
    .A2(_05497_),
    .B1(_05510_),
    .Y(_00871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_272 ();
 sky130_fd_sc_hd__nand2_1 _23451_ (.A(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .B(_05497_),
    .Y(_05512_));
 sky130_fd_sc_hd__o21ai_0 _23452_ (.A1(_02145_),
    .A2(_05497_),
    .B1(_05512_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_1 _23453_ (.A(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .B(_05497_),
    .Y(_05513_));
 sky130_fd_sc_hd__o21ai_0 _23454_ (.A1(_02297_),
    .A2(_05497_),
    .B1(_05513_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _23455_ (.A(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .B(_05497_),
    .Y(_05514_));
 sky130_fd_sc_hd__o21ai_0 _23456_ (.A1(_02414_),
    .A2(_05497_),
    .B1(_05514_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _23457_ (.A(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .B(_05497_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_0 _23458_ (.A1(_02535_),
    .A2(_05497_),
    .B1(_05515_),
    .Y(_00875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_271 ();
 sky130_fd_sc_hd__nand2_1 _23460_ (.A(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .B(_05497_),
    .Y(_05517_));
 sky130_fd_sc_hd__o21ai_0 _23461_ (.A1(_02628_),
    .A2(_05497_),
    .B1(_05517_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_1 _23462_ (.A(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .B(_05497_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21ai_0 _23463_ (.A1(net3453),
    .A2(_05497_),
    .B1(_05518_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _23464_ (.A(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .B(_05346_),
    .Y(_05519_));
 sky130_fd_sc_hd__o21ai_0 _23465_ (.A1(_02414_),
    .A2(_05346_),
    .B1(_05519_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _23466_ (.A(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .B(_05497_),
    .Y(_05520_));
 sky130_fd_sc_hd__o21ai_0 _23467_ (.A1(_02837_),
    .A2(_05497_),
    .B1(_05520_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _23468_ (.A(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .B(_05497_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_0 _23469_ (.A1(_02963_),
    .A2(_05497_),
    .B1(_05521_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_1 _23470_ (.A(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .B(_05497_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21ai_0 _23471_ (.A1(net3447),
    .A2(_05497_),
    .B1(_05522_),
    .Y(_00881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_270 ();
 sky130_fd_sc_hd__nor2_4 _23473_ (.A(_05147_),
    .B(_05466_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand2_1 _23474_ (.A(net3446),
    .B(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _23475_ (.A(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .B(_05497_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _23476_ (.A(_05525_),
    .B(_05526_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _23477_ (.A(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .B(_05497_),
    .Y(_05527_));
 sky130_fd_sc_hd__o21ai_0 _23478_ (.A1(net3425),
    .A2(_05497_),
    .B1(_05527_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _23479_ (.A(net3416),
    .B(_05524_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _23480_ (.A(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .B(_05497_),
    .Y(_05529_));
 sky130_fd_sc_hd__nand2_1 _23481_ (.A(_05528_),
    .B(_05529_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _23482_ (.A(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .B(_05497_),
    .Y(_05530_));
 sky130_fd_sc_hd__o21ai_0 _23483_ (.A1(net3433),
    .A2(_05497_),
    .B1(_05530_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _23484_ (.A(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .B(_05497_),
    .Y(_05531_));
 sky130_fd_sc_hd__o21ai_0 _23485_ (.A1(net3413),
    .A2(_05497_),
    .B1(_05531_),
    .Y(_00886_));
 sky130_fd_sc_hd__mux2_1 _23486_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A1(net3412),
    .S(_05524_),
    .X(_00887_));
 sky130_fd_sc_hd__nand2_1 _23487_ (.A(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .B(_05497_),
    .Y(_05532_));
 sky130_fd_sc_hd__o21ai_0 _23488_ (.A1(net3411),
    .A2(_05497_),
    .B1(_05532_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _23489_ (.A(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B(_05346_),
    .Y(_05533_));
 sky130_fd_sc_hd__o21ai_0 _23490_ (.A1(_02535_),
    .A2(_05346_),
    .B1(_05533_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand2_1 _23491_ (.A(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .B(_05497_),
    .Y(_05534_));
 sky130_fd_sc_hd__o21ai_0 _23492_ (.A1(net3410),
    .A2(_05497_),
    .B1(_05534_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _23493_ (.A(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .B(_05497_),
    .Y(_05535_));
 sky130_fd_sc_hd__o21ai_0 _23494_ (.A1(net3409),
    .A2(_05497_),
    .B1(_05535_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _23495_ (.A(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .B(_05497_),
    .Y(_05536_));
 sky130_fd_sc_hd__o21ai_0 _23496_ (.A1(net3408),
    .A2(_05497_),
    .B1(_05536_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand2_1 _23497_ (.A(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .B(_05497_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_0 _23498_ (.A1(net3407),
    .A2(_05497_),
    .B1(_05537_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand2_1 _23499_ (.A(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .B(_05497_),
    .Y(_05538_));
 sky130_fd_sc_hd__o21ai_0 _23500_ (.A1(net3406),
    .A2(_05497_),
    .B1(_05538_),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2_1 _23501_ (.A(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .B(_05524_),
    .Y(_05539_));
 sky130_fd_sc_hd__a31oi_1 _23502_ (.A1(net3405),
    .A2(net3457),
    .A3(_05524_),
    .B1(_05539_),
    .Y(_00895_));
 sky130_fd_sc_hd__mux2_1 _23503_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A1(net3404),
    .S(_05524_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_1 _23504_ (.A(_04920_),
    .B(_05497_),
    .Y(_05540_));
 sky130_fd_sc_hd__a22o_1 _23505_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .A2(_05497_),
    .B1(_05540_),
    .B2(net3403),
    .X(_00897_));
 sky130_fd_sc_hd__nand2_8 _23506_ (.A(_05165_),
    .B(_05428_),
    .Y(_05541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_267 ();
 sky130_fd_sc_hd__nand2_1 _23510_ (.A(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .B(_05541_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21ai_0 _23511_ (.A1(_05011_),
    .A2(_05541_),
    .B1(_05545_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2_1 _23512_ (.A(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .B(_05541_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_0 _23513_ (.A1(_05039_),
    .A2(_05541_),
    .B1(_05546_),
    .Y(_00899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_266 ();
 sky130_fd_sc_hd__nand2_1 _23515_ (.A(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .B(_05346_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_0 _23516_ (.A1(_02628_),
    .A2(_05346_),
    .B1(_05548_),
    .Y(_00900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_265 ();
 sky130_fd_sc_hd__nand2_1 _23518_ (.A(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .B(_05541_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_0 _23519_ (.A1(_05059_),
    .A2(_05541_),
    .B1(_05550_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _23520_ (.A(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .B(_05541_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21ai_0 _23521_ (.A1(net3463),
    .A2(_05541_),
    .B1(_05551_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_1 _23522_ (.A(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .B(_05541_),
    .Y(_05552_));
 sky130_fd_sc_hd__o21ai_0 _23523_ (.A1(net3459),
    .A2(_05541_),
    .B1(_05552_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_1 _23524_ (.A(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .B(_05541_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21ai_0 _23525_ (.A1(_04483_),
    .A2(_05541_),
    .B1(_05553_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _23526_ (.A(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .B(_05541_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_0 _23527_ (.A1(net3444),
    .A2(_05541_),
    .B1(_05554_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _23528_ (.A(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .B(_05541_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_0 _23529_ (.A1(_04964_),
    .A2(_05541_),
    .B1(_05555_),
    .Y(_00906_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_264 ();
 sky130_fd_sc_hd__nand2_1 _23531_ (.A(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .B(_05541_),
    .Y(_05557_));
 sky130_fd_sc_hd__o21ai_0 _23532_ (.A1(_02145_),
    .A2(_05541_),
    .B1(_05557_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand2_1 _23533_ (.A(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .B(_05541_),
    .Y(_05558_));
 sky130_fd_sc_hd__o21ai_0 _23534_ (.A1(_02297_),
    .A2(_05541_),
    .B1(_05558_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand2_1 _23535_ (.A(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .B(_05541_),
    .Y(_05559_));
 sky130_fd_sc_hd__o21ai_0 _23536_ (.A1(_02414_),
    .A2(_05541_),
    .B1(_05559_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_1 _23537_ (.A(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .B(_05541_),
    .Y(_05560_));
 sky130_fd_sc_hd__o21ai_0 _23538_ (.A1(_02535_),
    .A2(_05541_),
    .B1(_05560_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_1 _23539_ (.A(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .B(_05346_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_0 _23540_ (.A1(net3453),
    .A2(_05346_),
    .B1(_05561_),
    .Y(_00911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_263 ();
 sky130_fd_sc_hd__nand2_1 _23542_ (.A(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .B(_05541_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_0 _23543_ (.A1(_02628_),
    .A2(_05541_),
    .B1(_05563_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _23544_ (.A(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .B(_05541_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_0 _23545_ (.A1(net3453),
    .A2(_05541_),
    .B1(_05564_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _23546_ (.A(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .B(_05541_),
    .Y(_05565_));
 sky130_fd_sc_hd__o21ai_0 _23547_ (.A1(_02837_),
    .A2(_05541_),
    .B1(_05565_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _23548_ (.A(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .B(_05541_),
    .Y(_05566_));
 sky130_fd_sc_hd__o21ai_0 _23549_ (.A1(_02963_),
    .A2(_05541_),
    .B1(_05566_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_1 _23550_ (.A(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .B(_05541_),
    .Y(_05567_));
 sky130_fd_sc_hd__o21ai_0 _23551_ (.A1(net3447),
    .A2(_05541_),
    .B1(_05567_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_4 _23552_ (.A(_05191_),
    .B(_05466_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_1 _23553_ (.A(net3446),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _23554_ (.A(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .B(_05541_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_1 _23555_ (.A(_05569_),
    .B(_05570_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _23556_ (.A(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .B(_05541_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21ai_0 _23557_ (.A1(net3425),
    .A2(_05541_),
    .B1(_05571_),
    .Y(_00918_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_262 ();
 sky130_fd_sc_hd__nand2_1 _23559_ (.A(net3416),
    .B(_05568_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_1 _23560_ (.A(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .B(_05541_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_1 _23561_ (.A(_05573_),
    .B(_05574_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _23562_ (.A(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .B(_05541_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_0 _23563_ (.A1(net3433),
    .A2(_05541_),
    .B1(_05575_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_1 _23564_ (.A(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .B(_05541_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21ai_0 _23565_ (.A1(net3413),
    .A2(_05541_),
    .B1(_05576_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand2_1 _23566_ (.A(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .B(_05346_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_0 _23567_ (.A1(_02837_),
    .A2(_05346_),
    .B1(_05577_),
    .Y(_00922_));
 sky130_fd_sc_hd__mux2_1 _23568_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .A1(net3412),
    .S(_05568_),
    .X(_00923_));
 sky130_fd_sc_hd__nand2_1 _23569_ (.A(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .B(_05541_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21ai_0 _23570_ (.A1(net3411),
    .A2(_05541_),
    .B1(_05578_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _23571_ (.A(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .B(_05541_),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_0 _23572_ (.A1(net3410),
    .A2(_05541_),
    .B1(_05579_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _23573_ (.A(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .B(_05541_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_0 _23574_ (.A1(net3409),
    .A2(_05541_),
    .B1(_05580_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _23575_ (.A(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .B(_05541_),
    .Y(_05581_));
 sky130_fd_sc_hd__o21ai_0 _23576_ (.A1(net3408),
    .A2(_05541_),
    .B1(_05581_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_1 _23577_ (.A(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .B(_05541_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21ai_0 _23578_ (.A1(net3407),
    .A2(_05541_),
    .B1(_05582_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _23579_ (.A(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .B(_05541_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21ai_0 _23580_ (.A1(net3406),
    .A2(_05541_),
    .B1(_05583_),
    .Y(_00929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_260 ();
 sky130_fd_sc_hd__nor2_1 _23583_ (.A(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .B(_05568_),
    .Y(_05586_));
 sky130_fd_sc_hd__a31oi_1 _23584_ (.A1(net3405),
    .A2(net3457),
    .A3(_05568_),
    .B1(_05586_),
    .Y(_00930_));
 sky130_fd_sc_hd__mux2_1 _23585_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .A1(net3404),
    .S(_05568_),
    .X(_00931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_259 ();
 sky130_fd_sc_hd__nor2_1 _23587_ (.A(_04920_),
    .B(_05541_),
    .Y(_05588_));
 sky130_fd_sc_hd__a22o_1 _23588_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A2(_05541_),
    .B1(_05588_),
    .B2(net3403),
    .X(_00932_));
 sky130_fd_sc_hd__nand2_1 _23589_ (.A(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B(_05346_),
    .Y(_05589_));
 sky130_fd_sc_hd__o21ai_0 _23590_ (.A1(_02963_),
    .A2(_05346_),
    .B1(_05589_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_8 _23591_ (.A(_02151_),
    .B(_05428_),
    .Y(_05590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_256 ();
 sky130_fd_sc_hd__nand2_1 _23595_ (.A(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .B(_05590_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21ai_0 _23596_ (.A1(_05011_),
    .A2(_05590_),
    .B1(_05594_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_1 _23597_ (.A(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .B(_05590_),
    .Y(_05595_));
 sky130_fd_sc_hd__o21ai_0 _23598_ (.A1(net3456),
    .A2(_05590_),
    .B1(_05595_),
    .Y(_00935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_255 ();
 sky130_fd_sc_hd__nand2_1 _23600_ (.A(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .B(_05590_),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_0 _23601_ (.A1(_05059_),
    .A2(_05590_),
    .B1(_05597_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _23602_ (.A(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .B(_05590_),
    .Y(_05598_));
 sky130_fd_sc_hd__o21ai_0 _23603_ (.A1(net3463),
    .A2(_05590_),
    .B1(_05598_),
    .Y(_00937_));
 sky130_fd_sc_hd__nand2_1 _23604_ (.A(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .B(_05590_),
    .Y(_05599_));
 sky130_fd_sc_hd__o21ai_0 _23605_ (.A1(net3459),
    .A2(_05590_),
    .B1(_05599_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _23606_ (.A(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .B(_05590_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21ai_0 _23607_ (.A1(_04483_),
    .A2(_05590_),
    .B1(_05600_),
    .Y(_00939_));
 sky130_fd_sc_hd__nand2_1 _23608_ (.A(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .B(_05590_),
    .Y(_05601_));
 sky130_fd_sc_hd__o21ai_0 _23609_ (.A1(net3444),
    .A2(_05590_),
    .B1(_05601_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _23610_ (.A(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .B(_05590_),
    .Y(_05602_));
 sky130_fd_sc_hd__o21ai_0 _23611_ (.A1(_04964_),
    .A2(_05590_),
    .B1(_05602_),
    .Y(_00941_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_254 ();
 sky130_fd_sc_hd__nand2_1 _23613_ (.A(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .B(_05590_),
    .Y(_05604_));
 sky130_fd_sc_hd__o21ai_0 _23614_ (.A1(_02145_),
    .A2(_05590_),
    .B1(_05604_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand2_1 _23615_ (.A(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .B(_05590_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21ai_0 _23616_ (.A1(_02297_),
    .A2(_05590_),
    .B1(_05605_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _23617_ (.A(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .B(_05346_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _23618_ (.A1(net3447),
    .A2(_05346_),
    .B1(_05606_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand2_1 _23619_ (.A(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .B(_05590_),
    .Y(_05607_));
 sky130_fd_sc_hd__o21ai_0 _23620_ (.A1(_02414_),
    .A2(_05590_),
    .B1(_05607_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _23621_ (.A(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .B(_05590_),
    .Y(_05608_));
 sky130_fd_sc_hd__o21ai_0 _23622_ (.A1(_02535_),
    .A2(_05590_),
    .B1(_05608_),
    .Y(_00946_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_253 ();
 sky130_fd_sc_hd__nand2_1 _23624_ (.A(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .B(_05590_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21ai_0 _23625_ (.A1(_02628_),
    .A2(_05590_),
    .B1(_05610_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _23626_ (.A(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .B(_05590_),
    .Y(_05611_));
 sky130_fd_sc_hd__o21ai_0 _23627_ (.A1(net3453),
    .A2(_05590_),
    .B1(_05611_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _23628_ (.A(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .B(_05590_),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_0 _23629_ (.A1(_02837_),
    .A2(_05590_),
    .B1(_05612_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _23630_ (.A(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .B(_05590_),
    .Y(_05613_));
 sky130_fd_sc_hd__o21ai_0 _23631_ (.A1(_02963_),
    .A2(_05590_),
    .B1(_05613_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2_1 _23632_ (.A(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .B(_05590_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21ai_0 _23633_ (.A1(net3447),
    .A2(_05590_),
    .B1(_05614_),
    .Y(_00951_));
 sky130_fd_sc_hd__nor2_4 _23634_ (.A(_03094_),
    .B(_05466_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_1 _23635_ (.A(net3446),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _23636_ (.A(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .B(_05590_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand2_1 _23637_ (.A(_05616_),
    .B(_05617_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _23638_ (.A(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .B(_05590_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21ai_0 _23639_ (.A1(net3425),
    .A2(_05590_),
    .B1(_05618_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _23640_ (.A(net3416),
    .B(_05615_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand2_1 _23641_ (.A(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .B(_05590_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _23642_ (.A(_05619_),
    .B(_05620_),
    .Y(_00954_));
 sky130_fd_sc_hd__nor2_4 _23643_ (.A(_04978_),
    .B(_05147_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand2_1 _23644_ (.A(net3446),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _23645_ (.A(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .B(_05346_),
    .Y(_05623_));
 sky130_fd_sc_hd__nand2_1 _23646_ (.A(_05622_),
    .B(_05623_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _23647_ (.A(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .B(_05590_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_0 _23648_ (.A1(net3433),
    .A2(_05590_),
    .B1(_05624_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2_1 _23649_ (.A(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .B(_05590_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_0 _23650_ (.A1(net3413),
    .A2(_05590_),
    .B1(_05625_),
    .Y(_00957_));
 sky130_fd_sc_hd__mux2_1 _23651_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .A1(net3412),
    .S(_05615_),
    .X(_00958_));
 sky130_fd_sc_hd__nand2_1 _23652_ (.A(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .B(_05590_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_0 _23653_ (.A1(net3411),
    .A2(_05590_),
    .B1(_05626_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2_1 _23654_ (.A(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .B(_05590_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_0 _23655_ (.A1(net3410),
    .A2(_05590_),
    .B1(_05627_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _23656_ (.A(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .B(_05590_),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_0 _23657_ (.A1(net3409),
    .A2(_05590_),
    .B1(_05628_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_1 _23658_ (.A(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .B(_05590_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_0 _23659_ (.A1(net3408),
    .A2(_05590_),
    .B1(_05629_),
    .Y(_00962_));
 sky130_fd_sc_hd__nand2_1 _23660_ (.A(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .B(_05590_),
    .Y(_05630_));
 sky130_fd_sc_hd__o21ai_0 _23661_ (.A1(net3407),
    .A2(_05590_),
    .B1(_05630_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _23662_ (.A(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .B(_05590_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21ai_0 _23663_ (.A1(net3406),
    .A2(_05590_),
    .B1(_05631_),
    .Y(_00964_));
 sky130_fd_sc_hd__nor2_1 _23664_ (.A(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .B(_05615_),
    .Y(_05632_));
 sky130_fd_sc_hd__a31oi_1 _23665_ (.A1(net3405),
    .A2(net3457),
    .A3(_05615_),
    .B1(_05632_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _23666_ (.A(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B(_05346_),
    .Y(_05633_));
 sky130_fd_sc_hd__o21ai_0 _23667_ (.A1(net3425),
    .A2(_05346_),
    .B1(_05633_),
    .Y(_00966_));
 sky130_fd_sc_hd__mux2_1 _23668_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .A1(net3404),
    .S(_05615_),
    .X(_00967_));
 sky130_fd_sc_hd__nor2_1 _23669_ (.A(_04920_),
    .B(_05590_),
    .Y(_05634_));
 sky130_fd_sc_hd__a22o_1 _23670_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .A2(_05590_),
    .B1(_05634_),
    .B2(net3403),
    .X(_00968_));
 sky130_fd_sc_hd__nor2_4 _23671_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Y(_05635_));
 sky130_fd_sc_hd__and2_4 _23672_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .B(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__nand2_8 _23673_ (.A(_05015_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_250 ();
 sky130_fd_sc_hd__nand2_1 _23677_ (.A(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .B(_05637_),
    .Y(_05641_));
 sky130_fd_sc_hd__o21ai_0 _23678_ (.A1(_05011_),
    .A2(_05637_),
    .B1(_05641_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _23679_ (.A(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .B(_05637_),
    .Y(_05642_));
 sky130_fd_sc_hd__o21ai_0 _23680_ (.A1(net3456),
    .A2(_05637_),
    .B1(_05642_),
    .Y(_00970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_249 ();
 sky130_fd_sc_hd__nand2_1 _23682_ (.A(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .B(_05637_),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ai_0 _23683_ (.A1(_05059_),
    .A2(_05637_),
    .B1(_05644_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _23684_ (.A(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .B(_05637_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21ai_0 _23685_ (.A1(net3463),
    .A2(_05637_),
    .B1(_05645_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _23686_ (.A(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .B(_05637_),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ai_0 _23687_ (.A1(net3459),
    .A2(_05637_),
    .B1(_05646_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand2_1 _23688_ (.A(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .B(_05637_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_0 _23689_ (.A1(net3451),
    .A2(_05637_),
    .B1(_05647_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _23690_ (.A(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .B(_05637_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_0 _23691_ (.A1(net3444),
    .A2(_05637_),
    .B1(_05648_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _23692_ (.A(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .B(_05637_),
    .Y(_05649_));
 sky130_fd_sc_hd__o21ai_0 _23693_ (.A1(_04964_),
    .A2(_05637_),
    .B1(_05649_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _23694_ (.A(net3416),
    .B(_05621_),
    .Y(_05650_));
 sky130_fd_sc_hd__nand2_1 _23695_ (.A(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .B(_05346_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(_05650_),
    .B(_05651_),
    .Y(_00977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_248 ();
 sky130_fd_sc_hd__nand2_1 _23698_ (.A(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .B(_05637_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_0 _23699_ (.A1(_02145_),
    .A2(_05637_),
    .B1(_05653_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_1 _23700_ (.A(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .B(_05637_),
    .Y(_05654_));
 sky130_fd_sc_hd__o21ai_0 _23701_ (.A1(_02297_),
    .A2(_05637_),
    .B1(_05654_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _23702_ (.A(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .B(_05637_),
    .Y(_05655_));
 sky130_fd_sc_hd__o21ai_0 _23703_ (.A1(_02414_),
    .A2(_05637_),
    .B1(_05655_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _23704_ (.A(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .B(_05637_),
    .Y(_05656_));
 sky130_fd_sc_hd__o21ai_0 _23705_ (.A1(_02535_),
    .A2(_05637_),
    .B1(_05656_),
    .Y(_00981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_247 ();
 sky130_fd_sc_hd__nand2_1 _23707_ (.A(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .B(_05637_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_0 _23708_ (.A1(_02628_),
    .A2(_05637_),
    .B1(_05658_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _23709_ (.A(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .B(_05637_),
    .Y(_05659_));
 sky130_fd_sc_hd__o21ai_0 _23710_ (.A1(net3453),
    .A2(_05637_),
    .B1(_05659_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _23711_ (.A(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .B(_05637_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21ai_0 _23712_ (.A1(_02837_),
    .A2(_05637_),
    .B1(_05660_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _23713_ (.A(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .B(_05637_),
    .Y(_05661_));
 sky130_fd_sc_hd__o21ai_0 _23714_ (.A1(_02963_),
    .A2(_05637_),
    .B1(_05661_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _23715_ (.A(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .B(_05637_),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_0 _23716_ (.A1(net3447),
    .A2(_05637_),
    .B1(_05662_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_8 _23717_ (.A(net3945),
    .B(_05635_),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_4 _23718_ (.A(_05100_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _23719_ (.A(net3446),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__nand2_1 _23720_ (.A(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .B(_05637_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _23721_ (.A(_05665_),
    .B(_05666_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _23722_ (.A(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B(_05346_),
    .Y(_05667_));
 sky130_fd_sc_hd__o21ai_0 _23723_ (.A1(net3433),
    .A2(_05346_),
    .B1(_05667_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _23724_ (.A(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .B(_05637_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_0 _23725_ (.A1(net3425),
    .A2(_05637_),
    .B1(_05668_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _23726_ (.A(net3416),
    .B(_05664_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_1 _23727_ (.A(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .B(_05637_),
    .Y(_05670_));
 sky130_fd_sc_hd__nand2_1 _23728_ (.A(_05669_),
    .B(_05670_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand2_1 _23729_ (.A(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .B(_05637_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21ai_0 _23730_ (.A1(net3433),
    .A2(_05637_),
    .B1(_05671_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_1 _23731_ (.A(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .B(_05637_),
    .Y(_05672_));
 sky130_fd_sc_hd__o21ai_0 _23732_ (.A1(net3413),
    .A2(_05637_),
    .B1(_05672_),
    .Y(_00992_));
 sky130_fd_sc_hd__mux2_1 _23733_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A1(net3412),
    .S(_05664_),
    .X(_00993_));
 sky130_fd_sc_hd__nand2_1 _23734_ (.A(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .B(_05637_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21ai_0 _23735_ (.A1(net3411),
    .A2(_05637_),
    .B1(_05673_),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_1 _23736_ (.A(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .B(_05637_),
    .Y(_05674_));
 sky130_fd_sc_hd__o21ai_0 _23737_ (.A1(net3410),
    .A2(_05637_),
    .B1(_05674_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _23738_ (.A(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .B(_05637_),
    .Y(_05675_));
 sky130_fd_sc_hd__o21ai_0 _23739_ (.A1(net3409),
    .A2(_05637_),
    .B1(_05675_),
    .Y(_00996_));
 sky130_fd_sc_hd__nand2_1 _23740_ (.A(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .B(_05637_),
    .Y(_05676_));
 sky130_fd_sc_hd__o21ai_0 _23741_ (.A1(net3408),
    .A2(_05637_),
    .B1(_05676_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _23742_ (.A(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .B(_05637_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21ai_0 _23743_ (.A1(net3407),
    .A2(_05637_),
    .B1(_05677_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _23744_ (.A(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .B(_05346_),
    .Y(_05678_));
 sky130_fd_sc_hd__o21ai_0 _23745_ (.A1(net3413),
    .A2(_05346_),
    .B1(_05678_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _23746_ (.A(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .B(_05637_),
    .Y(_05679_));
 sky130_fd_sc_hd__o21ai_0 _23747_ (.A1(net3406),
    .A2(_05637_),
    .B1(_05679_),
    .Y(_01000_));
 sky130_fd_sc_hd__nor2_1 _23748_ (.A(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .B(_05664_),
    .Y(_05680_));
 sky130_fd_sc_hd__a31oi_1 _23749_ (.A1(net3405),
    .A2(net3457),
    .A3(_05664_),
    .B1(_05680_),
    .Y(_01001_));
 sky130_fd_sc_hd__mux2_1 _23750_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A1(net3404),
    .S(_05664_),
    .X(_01002_));
 sky130_fd_sc_hd__nor2_1 _23751_ (.A(net3464),
    .B(_05637_),
    .Y(_05681_));
 sky130_fd_sc_hd__a22o_1 _23752_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A2(_05637_),
    .B1(_05681_),
    .B2(net3403),
    .X(_01003_));
 sky130_fd_sc_hd__nand2_8 _23753_ (.A(_05122_),
    .B(_05636_),
    .Y(_05682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_244 ();
 sky130_fd_sc_hd__nand2_1 _23757_ (.A(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .B(_05682_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_0 _23758_ (.A1(_05011_),
    .A2(_05682_),
    .B1(_05686_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand2_1 _23759_ (.A(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .B(_05682_),
    .Y(_05687_));
 sky130_fd_sc_hd__o21ai_0 _23760_ (.A1(net3456),
    .A2(_05682_),
    .B1(_05687_),
    .Y(_01005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_243 ();
 sky130_fd_sc_hd__nand2_1 _23762_ (.A(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .B(_05682_),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ai_0 _23763_ (.A1(_05059_),
    .A2(_05682_),
    .B1(_05689_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_1 _23764_ (.A(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .B(_05682_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_0 _23765_ (.A1(net3463),
    .A2(_05682_),
    .B1(_05690_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _23766_ (.A(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .B(_05682_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21ai_0 _23767_ (.A1(net3459),
    .A2(_05682_),
    .B1(_05691_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_1 _23768_ (.A(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .B(_05682_),
    .Y(_05692_));
 sky130_fd_sc_hd__o21ai_0 _23769_ (.A1(net3451),
    .A2(_05682_),
    .B1(_05692_),
    .Y(_01009_));
 sky130_fd_sc_hd__mux2_1 _23770_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A1(net3412),
    .S(_05621_),
    .X(_01010_));
 sky130_fd_sc_hd__nand2_1 _23771_ (.A(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .B(_05682_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_0 _23772_ (.A1(net3444),
    .A2(_05682_),
    .B1(_05693_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _23773_ (.A(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .B(_05682_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_0 _23774_ (.A1(_04964_),
    .A2(_05682_),
    .B1(_05694_),
    .Y(_01012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_242 ();
 sky130_fd_sc_hd__nand2_1 _23776_ (.A(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .B(_05682_),
    .Y(_05696_));
 sky130_fd_sc_hd__o21ai_0 _23777_ (.A1(_02145_),
    .A2(_05682_),
    .B1(_05696_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _23778_ (.A(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .B(_05682_),
    .Y(_05697_));
 sky130_fd_sc_hd__o21ai_0 _23779_ (.A1(_02297_),
    .A2(_05682_),
    .B1(_05697_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _23780_ (.A(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .B(_05682_),
    .Y(_05698_));
 sky130_fd_sc_hd__o21ai_0 _23781_ (.A1(_02414_),
    .A2(_05682_),
    .B1(_05698_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _23782_ (.A(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .B(_05682_),
    .Y(_05699_));
 sky130_fd_sc_hd__o21ai_0 _23783_ (.A1(_02535_),
    .A2(_05682_),
    .B1(_05699_),
    .Y(_01016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_241 ();
 sky130_fd_sc_hd__nand2_1 _23785_ (.A(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .B(_05682_),
    .Y(_05701_));
 sky130_fd_sc_hd__o21ai_0 _23786_ (.A1(_02628_),
    .A2(_05682_),
    .B1(_05701_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _23787_ (.A(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .B(_05682_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_0 _23788_ (.A1(net3453),
    .A2(_05682_),
    .B1(_05702_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _23789_ (.A(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .B(_05682_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_0 _23790_ (.A1(_02837_),
    .A2(_05682_),
    .B1(_05703_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _23791_ (.A(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .B(_05682_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_0 _23792_ (.A1(_02963_),
    .A2(_05682_),
    .B1(_05704_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _23793_ (.A(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .B(_05346_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_0 _23794_ (.A1(net3411),
    .A2(_05346_),
    .B1(_05705_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _23795_ (.A(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .B(_05682_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_0 _23796_ (.A1(net3447),
    .A2(_05682_),
    .B1(_05706_),
    .Y(_01022_));
 sky130_fd_sc_hd__nor2_4 _23797_ (.A(_05147_),
    .B(_05663_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_1 _23798_ (.A(net3446),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _23799_ (.A(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .B(_05682_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_1 _23800_ (.A(_05708_),
    .B(_05709_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_1 _23801_ (.A(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .B(_05682_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21ai_0 _23802_ (.A1(net3425),
    .A2(_05682_),
    .B1(_05710_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _23803_ (.A(net3416),
    .B(_05707_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2_1 _23804_ (.A(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .B(_05682_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _23805_ (.A(_05711_),
    .B(_05712_),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2_1 _23806_ (.A(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .B(_05682_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _23807_ (.A1(net3433),
    .A2(_05682_),
    .B1(_05713_),
    .Y(_01026_));
 sky130_fd_sc_hd__nand2_1 _23808_ (.A(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .B(_05682_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_0 _23809_ (.A1(net3413),
    .A2(_05682_),
    .B1(_05714_),
    .Y(_01027_));
 sky130_fd_sc_hd__mux2_1 _23810_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A1(net3412),
    .S(_05707_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_1 _23811_ (.A(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .B(_05682_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ai_0 _23812_ (.A1(net3411),
    .A2(_05682_),
    .B1(_05715_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _23813_ (.A(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .B(_05682_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_0 _23814_ (.A1(net3410),
    .A2(_05682_),
    .B1(_05716_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_1 _23815_ (.A(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .B(_05682_),
    .Y(_05717_));
 sky130_fd_sc_hd__o21ai_0 _23816_ (.A1(net3409),
    .A2(_05682_),
    .B1(_05717_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _23817_ (.A(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .B(_05346_),
    .Y(_05718_));
 sky130_fd_sc_hd__o21ai_0 _23818_ (.A1(net3410),
    .A2(_05346_),
    .B1(_05718_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _23819_ (.A(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .B(_05682_),
    .Y(_05719_));
 sky130_fd_sc_hd__o21ai_0 _23820_ (.A1(net3408),
    .A2(_05682_),
    .B1(_05719_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _23821_ (.A(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .B(_05682_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_0 _23822_ (.A1(net3407),
    .A2(_05682_),
    .B1(_05720_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _23823_ (.A(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .B(_05682_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21ai_0 _23824_ (.A1(net3406),
    .A2(_05682_),
    .B1(_05721_),
    .Y(_01035_));
 sky130_fd_sc_hd__nor2_1 _23825_ (.A(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .B(_05707_),
    .Y(_05722_));
 sky130_fd_sc_hd__a31oi_1 _23826_ (.A1(net3405),
    .A2(net3457),
    .A3(_05707_),
    .B1(_05722_),
    .Y(_01036_));
 sky130_fd_sc_hd__mux2_1 _23827_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .A1(net3404),
    .S(_05707_),
    .X(_01037_));
 sky130_fd_sc_hd__nor2_1 _23828_ (.A(net3464),
    .B(_05682_),
    .Y(_05723_));
 sky130_fd_sc_hd__a22o_1 _23829_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A2(_05682_),
    .B1(_05723_),
    .B2(net3403),
    .X(_01038_));
 sky130_fd_sc_hd__nand2_8 _23830_ (.A(_05165_),
    .B(_05636_),
    .Y(_05724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_238 ();
 sky130_fd_sc_hd__nand2_1 _23834_ (.A(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .B(_05724_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_0 _23835_ (.A1(_05011_),
    .A2(_05724_),
    .B1(_05728_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_1 _23836_ (.A(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .B(_05724_),
    .Y(_05729_));
 sky130_fd_sc_hd__o21ai_0 _23837_ (.A1(net3456),
    .A2(_05724_),
    .B1(_05729_),
    .Y(_01040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_237 ();
 sky130_fd_sc_hd__nand2_1 _23839_ (.A(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .B(_05724_),
    .Y(_05731_));
 sky130_fd_sc_hd__o21ai_0 _23840_ (.A1(_05059_),
    .A2(_05724_),
    .B1(_05731_),
    .Y(_01041_));
 sky130_fd_sc_hd__nand2_1 _23841_ (.A(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .B(_05724_),
    .Y(_05732_));
 sky130_fd_sc_hd__o21ai_0 _23842_ (.A1(net3463),
    .A2(_05724_),
    .B1(_05732_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _23843_ (.A(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .B(_05346_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_0 _23844_ (.A1(net3409),
    .A2(_05346_),
    .B1(_05733_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _23845_ (.A(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .B(_05724_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21ai_0 _23846_ (.A1(net3459),
    .A2(_05724_),
    .B1(_05734_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand2_1 _23847_ (.A(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .B(_05724_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_0 _23848_ (.A1(net3451),
    .A2(_05724_),
    .B1(_05735_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand2_1 _23849_ (.A(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .B(_05724_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_0 _23850_ (.A1(net3444),
    .A2(_05724_),
    .B1(_05736_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _23851_ (.A(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .B(_05724_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21ai_0 _23852_ (.A1(_04964_),
    .A2(_05724_),
    .B1(_05737_),
    .Y(_01047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_236 ();
 sky130_fd_sc_hd__nand2_1 _23854_ (.A(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .B(_05724_),
    .Y(_05739_));
 sky130_fd_sc_hd__o21ai_0 _23855_ (.A1(_02145_),
    .A2(_05724_),
    .B1(_05739_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand2_1 _23856_ (.A(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .B(_05724_),
    .Y(_05740_));
 sky130_fd_sc_hd__o21ai_0 _23857_ (.A1(_02297_),
    .A2(_05724_),
    .B1(_05740_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _23858_ (.A(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .B(_05724_),
    .Y(_05741_));
 sky130_fd_sc_hd__o21ai_0 _23859_ (.A1(_02414_),
    .A2(_05724_),
    .B1(_05741_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _23860_ (.A(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .B(_05724_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21ai_0 _23861_ (.A1(_02535_),
    .A2(_05724_),
    .B1(_05742_),
    .Y(_01051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_235 ();
 sky130_fd_sc_hd__nand2_1 _23863_ (.A(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .B(_05724_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_0 _23864_ (.A1(_02628_),
    .A2(_05724_),
    .B1(_05744_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _23865_ (.A(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .B(_05724_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_0 _23866_ (.A1(net3453),
    .A2(_05724_),
    .B1(_05745_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand2_1 _23867_ (.A(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B(_05346_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _23868_ (.A1(net3408),
    .A2(_05346_),
    .B1(_05746_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _23869_ (.A(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .B(_05724_),
    .Y(_05747_));
 sky130_fd_sc_hd__o21ai_0 _23870_ (.A1(_02837_),
    .A2(_05724_),
    .B1(_05747_),
    .Y(_01055_));
 sky130_fd_sc_hd__nand2_1 _23871_ (.A(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .B(_05724_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_0 _23872_ (.A1(_02963_),
    .A2(_05724_),
    .B1(_05748_),
    .Y(_01056_));
 sky130_fd_sc_hd__nand2_1 _23873_ (.A(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .B(_05724_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_0 _23874_ (.A1(net3447),
    .A2(_05724_),
    .B1(_05749_),
    .Y(_01057_));
 sky130_fd_sc_hd__nor2_4 _23875_ (.A(_05191_),
    .B(_05663_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_1 _23876_ (.A(net3446),
    .B(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand2_1 _23877_ (.A(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .B(_05724_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_1 _23878_ (.A(_05751_),
    .B(_05752_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_1 _23879_ (.A(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .B(_05724_),
    .Y(_05753_));
 sky130_fd_sc_hd__o21ai_0 _23880_ (.A1(net3425),
    .A2(_05724_),
    .B1(_05753_),
    .Y(_01059_));
 sky130_fd_sc_hd__nand2_1 _23881_ (.A(net3416),
    .B(_05750_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _23882_ (.A(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .B(_05724_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _23883_ (.A(_05754_),
    .B(_05755_),
    .Y(_01060_));
 sky130_fd_sc_hd__nand2_1 _23884_ (.A(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .B(_05724_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_0 _23885_ (.A1(net3433),
    .A2(_05724_),
    .B1(_05756_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand2_1 _23886_ (.A(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .B(_05724_),
    .Y(_05757_));
 sky130_fd_sc_hd__o21ai_0 _23887_ (.A1(net3413),
    .A2(_05724_),
    .B1(_05757_),
    .Y(_01062_));
 sky130_fd_sc_hd__mux2_1 _23888_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .A1(net3412),
    .S(_05750_),
    .X(_01063_));
 sky130_fd_sc_hd__nand2_1 _23889_ (.A(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .B(_05724_),
    .Y(_05758_));
 sky130_fd_sc_hd__o21ai_0 _23890_ (.A1(net3411),
    .A2(_05724_),
    .B1(_05758_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _23891_ (.A(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .B(_05346_),
    .Y(_05759_));
 sky130_fd_sc_hd__o21ai_0 _23892_ (.A1(net3407),
    .A2(_05346_),
    .B1(_05759_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand2_1 _23893_ (.A(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .B(_05724_),
    .Y(_05760_));
 sky130_fd_sc_hd__o21ai_0 _23894_ (.A1(net3410),
    .A2(_05724_),
    .B1(_05760_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _23895_ (.A(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .B(_05724_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_0 _23896_ (.A1(net3409),
    .A2(_05724_),
    .B1(_05761_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _23897_ (.A(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .B(_05724_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_0 _23898_ (.A1(net3408),
    .A2(_05724_),
    .B1(_05762_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _23899_ (.A(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .B(_05724_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21ai_0 _23900_ (.A1(net3407),
    .A2(_05724_),
    .B1(_05763_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _23901_ (.A(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .B(_05724_),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_0 _23902_ (.A1(net3406),
    .A2(_05724_),
    .B1(_05764_),
    .Y(_01070_));
 sky130_fd_sc_hd__nor2_1 _23903_ (.A(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .B(_05750_),
    .Y(_05765_));
 sky130_fd_sc_hd__a31oi_1 _23904_ (.A1(net3405),
    .A2(net3457),
    .A3(_05750_),
    .B1(_05765_),
    .Y(_01071_));
 sky130_fd_sc_hd__mux2_1 _23905_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .A1(net3404),
    .S(_05750_),
    .X(_01072_));
 sky130_fd_sc_hd__nor2_1 _23906_ (.A(net3464),
    .B(_05724_),
    .Y(_05766_));
 sky130_fd_sc_hd__a22o_1 _23907_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A2(_05724_),
    .B1(_05766_),
    .B2(net3403),
    .X(_01073_));
 sky130_fd_sc_hd__nand2_8 _23908_ (.A(_02151_),
    .B(_05636_),
    .Y(_05767_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_232 ();
 sky130_fd_sc_hd__nand2_1 _23912_ (.A(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .B(_05767_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_0 _23913_ (.A1(_05011_),
    .A2(_05767_),
    .B1(_05771_),
    .Y(_01074_));
 sky130_fd_sc_hd__nand2_1 _23914_ (.A(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .B(_05767_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_0 _23915_ (.A1(net3456),
    .A2(_05767_),
    .B1(_05772_),
    .Y(_01075_));
 sky130_fd_sc_hd__nand2_1 _23916_ (.A(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .B(_05346_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21ai_0 _23917_ (.A1(net3406),
    .A2(_05346_),
    .B1(_05773_),
    .Y(_01076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 ();
 sky130_fd_sc_hd__nand2_1 _23919_ (.A(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .B(_05767_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ai_0 _23920_ (.A1(_05059_),
    .A2(_05767_),
    .B1(_05775_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand2_1 _23921_ (.A(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .B(_05767_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_0 _23922_ (.A1(net3463),
    .A2(_05767_),
    .B1(_05776_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _23923_ (.A(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .B(_05767_),
    .Y(_05777_));
 sky130_fd_sc_hd__o21ai_0 _23924_ (.A1(net3459),
    .A2(_05767_),
    .B1(_05777_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2_1 _23925_ (.A(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .B(_05767_),
    .Y(_05778_));
 sky130_fd_sc_hd__o21ai_0 _23926_ (.A1(net3451),
    .A2(_05767_),
    .B1(_05778_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _23927_ (.A(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .B(_05767_),
    .Y(_05779_));
 sky130_fd_sc_hd__o21ai_0 _23928_ (.A1(net3444),
    .A2(_05767_),
    .B1(_05779_),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _23929_ (.A(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .B(_05767_),
    .Y(_05780_));
 sky130_fd_sc_hd__o21ai_0 _23930_ (.A1(_04964_),
    .A2(_05767_),
    .B1(_05780_),
    .Y(_01082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 ();
 sky130_fd_sc_hd__nand2_1 _23932_ (.A(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .B(_05767_),
    .Y(_05782_));
 sky130_fd_sc_hd__o21ai_0 _23933_ (.A1(_02145_),
    .A2(_05767_),
    .B1(_05782_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _23934_ (.A(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .B(_05767_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_0 _23935_ (.A1(_02297_),
    .A2(_05767_),
    .B1(_05783_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand2_1 _23936_ (.A(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .B(_05767_),
    .Y(_05784_));
 sky130_fd_sc_hd__o21ai_0 _23937_ (.A1(_02414_),
    .A2(_05767_),
    .B1(_05784_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _23938_ (.A(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .B(_05767_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ai_0 _23939_ (.A1(_02535_),
    .A2(_05767_),
    .B1(_05785_),
    .Y(_01086_));
 sky130_fd_sc_hd__nor2_1 _23940_ (.A(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .B(_05621_),
    .Y(_05786_));
 sky130_fd_sc_hd__a31oi_1 _23941_ (.A1(net3405),
    .A2(net3457),
    .A3(_05621_),
    .B1(_05786_),
    .Y(_01087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 ();
 sky130_fd_sc_hd__nand2_1 _23943_ (.A(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .B(_05767_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_0 _23944_ (.A1(_02628_),
    .A2(_05767_),
    .B1(_05788_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _23945_ (.A(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .B(_05767_),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_0 _23946_ (.A1(net3453),
    .A2(_05767_),
    .B1(_05789_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _23947_ (.A(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .B(_05767_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_0 _23948_ (.A1(_02837_),
    .A2(_05767_),
    .B1(_05790_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _23949_ (.A(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .B(_05767_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_0 _23950_ (.A1(_02963_),
    .A2(_05767_),
    .B1(_05791_),
    .Y(_01091_));
 sky130_fd_sc_hd__nand2_1 _23951_ (.A(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .B(_05767_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ai_0 _23952_ (.A1(net3447),
    .A2(_05767_),
    .B1(_05792_),
    .Y(_01092_));
 sky130_fd_sc_hd__nor2_4 _23953_ (.A(_03094_),
    .B(_05663_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _23954_ (.A(net3446),
    .B(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__nand2_1 _23955_ (.A(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .B(_05767_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(_05794_),
    .B(_05795_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand2_1 _23957_ (.A(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .B(_05767_),
    .Y(_05796_));
 sky130_fd_sc_hd__o21ai_0 _23958_ (.A1(net3425),
    .A2(_05767_),
    .B1(_05796_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand2_1 _23959_ (.A(net3416),
    .B(_05793_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_1 _23960_ (.A(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .B(_05767_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _23961_ (.A(_05797_),
    .B(_05798_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand2_1 _23962_ (.A(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .B(_05767_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_0 _23963_ (.A1(net3433),
    .A2(_05767_),
    .B1(_05799_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _23964_ (.A(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .B(_05767_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_0 _23965_ (.A1(net3413),
    .A2(_05767_),
    .B1(_05800_),
    .Y(_01097_));
 sky130_fd_sc_hd__mux2_1 _23966_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A1(net3404),
    .S(_05621_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _23967_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .A1(net3412),
    .S(_05793_),
    .X(_01099_));
 sky130_fd_sc_hd__nand2_1 _23968_ (.A(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .B(_05767_),
    .Y(_05801_));
 sky130_fd_sc_hd__o21ai_0 _23969_ (.A1(net3411),
    .A2(_05767_),
    .B1(_05801_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _23970_ (.A(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .B(_05767_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_0 _23971_ (.A1(net3410),
    .A2(_05767_),
    .B1(_05802_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _23972_ (.A(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .B(_05767_),
    .Y(_05803_));
 sky130_fd_sc_hd__o21ai_0 _23973_ (.A1(net3409),
    .A2(_05767_),
    .B1(_05803_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _23974_ (.A(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .B(_05767_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_0 _23975_ (.A1(net3408),
    .A2(_05767_),
    .B1(_05804_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _23976_ (.A(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .B(_05767_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _23977_ (.A1(net3407),
    .A2(_05767_),
    .B1(_05805_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _23978_ (.A(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .B(_05767_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_0 _23979_ (.A1(net3406),
    .A2(_05767_),
    .B1(_05806_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _23980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .B(_05793_),
    .Y(_05807_));
 sky130_fd_sc_hd__a31oi_1 _23981_ (.A1(net3405),
    .A2(net3457),
    .A3(_05793_),
    .B1(_05807_),
    .Y(_01106_));
 sky130_fd_sc_hd__mux2_1 _23982_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .A1(net3404),
    .S(_05793_),
    .X(_01107_));
 sky130_fd_sc_hd__nor2_1 _23983_ (.A(net3464),
    .B(_05767_),
    .Y(_05808_));
 sky130_fd_sc_hd__a22o_1 _23984_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .A2(_05767_),
    .B1(_05808_),
    .B2(net3403),
    .X(_01108_));
 sky130_fd_sc_hd__nor2_1 _23985_ (.A(_04920_),
    .B(_05346_),
    .Y(_05809_));
 sky130_fd_sc_hd__a22o_1 _23986_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A2(_05346_),
    .B1(_05809_),
    .B2(net3403),
    .X(_01109_));
 sky130_fd_sc_hd__and3b_4 _23987_ (.A_N(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .X(_05810_));
 sky130_fd_sc_hd__nand2_8 _23988_ (.A(_05015_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__nand2_1 _23992_ (.A(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .B(_05811_),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_0 _23993_ (.A1(_05011_),
    .A2(_05811_),
    .B1(_05815_),
    .Y(_01110_));
 sky130_fd_sc_hd__nand2_1 _23994_ (.A(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .B(_05811_),
    .Y(_05816_));
 sky130_fd_sc_hd__o21ai_0 _23995_ (.A1(net3456),
    .A2(_05811_),
    .B1(_05816_),
    .Y(_01111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__nand2_1 _23997_ (.A(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .B(_05811_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_0 _23998_ (.A1(_05059_),
    .A2(_05811_),
    .B1(_05818_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _23999_ (.A(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .B(_05811_),
    .Y(_05819_));
 sky130_fd_sc_hd__o21ai_0 _24000_ (.A1(net3463),
    .A2(_05811_),
    .B1(_05819_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _24001_ (.A(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .B(_05811_),
    .Y(_05820_));
 sky130_fd_sc_hd__o21ai_0 _24002_ (.A1(net3459),
    .A2(_05811_),
    .B1(_05820_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2_1 _24003_ (.A(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .B(_05811_),
    .Y(_05821_));
 sky130_fd_sc_hd__o21ai_0 _24004_ (.A1(net3451),
    .A2(_05811_),
    .B1(_05821_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _24005_ (.A(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .B(_05811_),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_0 _24006_ (.A1(net3444),
    .A2(_05811_),
    .B1(_05822_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _24007_ (.A(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .B(_05811_),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_0 _24008_ (.A1(_04964_),
    .A2(_05811_),
    .B1(_05823_),
    .Y(_01117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__nand2_1 _24010_ (.A(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .B(_05811_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ai_0 _24011_ (.A1(_02145_),
    .A2(_05811_),
    .B1(_05825_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_1 _24012_ (.A(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .B(_05811_),
    .Y(_05826_));
 sky130_fd_sc_hd__o21ai_0 _24013_ (.A1(_02297_),
    .A2(_05811_),
    .B1(_05826_),
    .Y(_01119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__nand2_8 _24015_ (.A(_10519_),
    .B(_05165_),
    .Y(_05828_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_220 ();
 sky130_fd_sc_hd__nand2_1 _24019_ (.A(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .B(_05828_),
    .Y(_05832_));
 sky130_fd_sc_hd__o21ai_0 _24020_ (.A1(_05011_),
    .A2(_05828_),
    .B1(_05832_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _24021_ (.A(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .B(_05811_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_0 _24022_ (.A1(_02414_),
    .A2(_05811_),
    .B1(_05833_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _24023_ (.A(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .B(_05811_),
    .Y(_05834_));
 sky130_fd_sc_hd__o21ai_0 _24024_ (.A1(_02535_),
    .A2(_05811_),
    .B1(_05834_),
    .Y(_01122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_219 ();
 sky130_fd_sc_hd__nand2_1 _24026_ (.A(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .B(_05811_),
    .Y(_05836_));
 sky130_fd_sc_hd__o21ai_0 _24027_ (.A1(_02628_),
    .A2(_05811_),
    .B1(_05836_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand2_1 _24028_ (.A(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .B(_05811_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_0 _24029_ (.A1(net3453),
    .A2(_05811_),
    .B1(_05837_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _24030_ (.A(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .B(_05811_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ai_0 _24031_ (.A1(_02837_),
    .A2(_05811_),
    .B1(_05838_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _24032_ (.A(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .B(_05811_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_0 _24033_ (.A1(_02963_),
    .A2(_05811_),
    .B1(_05839_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand2_1 _24034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .B(_05811_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21ai_0 _24035_ (.A1(net3447),
    .A2(_05811_),
    .B1(_05840_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand3b_1 _24036_ (.A_N(net3946),
    .B(net3827),
    .C(net3945),
    .Y(_05841_));
 sky130_fd_sc_hd__nor2_4 _24037_ (.A(_05100_),
    .B(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand2_1 _24038_ (.A(net3446),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_1 _24039_ (.A(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .B(_05811_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_1 _24040_ (.A(_05843_),
    .B(_05844_),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _24041_ (.A(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .B(_05811_),
    .Y(_05845_));
 sky130_fd_sc_hd__o21ai_0 _24042_ (.A1(net3425),
    .A2(_05811_),
    .B1(_05845_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _24043_ (.A(net3416),
    .B(_05842_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _24044_ (.A(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .B(_05811_),
    .Y(_05847_));
 sky130_fd_sc_hd__nand2_1 _24045_ (.A(_05846_),
    .B(_05847_),
    .Y(_01130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_218 ();
 sky130_fd_sc_hd__nand2_1 _24047_ (.A(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .B(_05828_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21ai_0 _24048_ (.A1(_05039_),
    .A2(_05828_),
    .B1(_05849_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _24049_ (.A(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .B(_05811_),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_0 _24050_ (.A1(net3433),
    .A2(_05811_),
    .B1(_05850_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _24051_ (.A(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .B(_05811_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_0 _24052_ (.A1(net3413),
    .A2(_05811_),
    .B1(_05851_),
    .Y(_01133_));
 sky130_fd_sc_hd__mux2_1 _24053_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(net3412),
    .S(_05842_),
    .X(_01134_));
 sky130_fd_sc_hd__nand2_1 _24054_ (.A(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .B(_05811_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_0 _24055_ (.A1(net3411),
    .A2(_05811_),
    .B1(_05852_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _24056_ (.A(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .B(_05811_),
    .Y(_05853_));
 sky130_fd_sc_hd__o21ai_0 _24057_ (.A1(net3410),
    .A2(_05811_),
    .B1(_05853_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand2_1 _24058_ (.A(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .B(_05811_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_0 _24059_ (.A1(net3409),
    .A2(_05811_),
    .B1(_05854_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2_1 _24060_ (.A(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .B(_05811_),
    .Y(_05855_));
 sky130_fd_sc_hd__o21ai_0 _24061_ (.A1(net3408),
    .A2(_05811_),
    .B1(_05855_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2_1 _24062_ (.A(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .B(_05811_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _24063_ (.A1(net3407),
    .A2(_05811_),
    .B1(_05856_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _24064_ (.A(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .B(_05811_),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_0 _24065_ (.A1(net3406),
    .A2(_05811_),
    .B1(_05857_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _24066_ (.A(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .B(_05842_),
    .Y(_05858_));
 sky130_fd_sc_hd__a31oi_1 _24067_ (.A1(net3405),
    .A2(net3457),
    .A3(_05842_),
    .B1(_05858_),
    .Y(_01141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_216 ();
 sky130_fd_sc_hd__nand2_1 _24070_ (.A(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .B(_05828_),
    .Y(_05861_));
 sky130_fd_sc_hd__o21ai_0 _24071_ (.A1(_05059_),
    .A2(_05828_),
    .B1(_05861_),
    .Y(_01142_));
 sky130_fd_sc_hd__mux2_1 _24072_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A1(net3404),
    .S(_05842_),
    .X(_01143_));
 sky130_fd_sc_hd__nor2_1 _24073_ (.A(net3464),
    .B(_05811_),
    .Y(_05862_));
 sky130_fd_sc_hd__a22o_1 _24074_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A2(_05811_),
    .B1(_05862_),
    .B2(net3403),
    .X(_01144_));
 sky130_fd_sc_hd__nand2_8 _24075_ (.A(_05122_),
    .B(_05810_),
    .Y(_05863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_213 ();
 sky130_fd_sc_hd__nand2_1 _24079_ (.A(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .B(_05863_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_0 _24080_ (.A1(_05011_),
    .A2(_05863_),
    .B1(_05867_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .B(_05863_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_0 _24082_ (.A1(net3456),
    .A2(_05863_),
    .B1(_05868_),
    .Y(_01146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_212 ();
 sky130_fd_sc_hd__nand2_1 _24084_ (.A(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .B(_05863_),
    .Y(_05870_));
 sky130_fd_sc_hd__o21ai_0 _24085_ (.A1(_05059_),
    .A2(_05863_),
    .B1(_05870_),
    .Y(_01147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_211 ();
 sky130_fd_sc_hd__nand2_1 _24087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .B(_05863_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_0 _24088_ (.A1(net3463),
    .A2(_05863_),
    .B1(_05872_),
    .Y(_01148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_210 ();
 sky130_fd_sc_hd__nand2_1 _24090_ (.A(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .B(_05863_),
    .Y(_05874_));
 sky130_fd_sc_hd__o21ai_0 _24091_ (.A1(net3459),
    .A2(_05863_),
    .B1(_05874_),
    .Y(_01149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_209 ();
 sky130_fd_sc_hd__nand2_1 _24093_ (.A(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .B(_05863_),
    .Y(_05876_));
 sky130_fd_sc_hd__o21ai_0 _24094_ (.A1(net3451),
    .A2(_05863_),
    .B1(_05876_),
    .Y(_01150_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_208 ();
 sky130_fd_sc_hd__nand2_1 _24096_ (.A(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .B(_05863_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21ai_0 _24097_ (.A1(net3444),
    .A2(_05863_),
    .B1(_05878_),
    .Y(_01151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_207 ();
 sky130_fd_sc_hd__nand2_1 _24099_ (.A(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .B(_05863_),
    .Y(_05880_));
 sky130_fd_sc_hd__o21ai_0 _24100_ (.A1(_04964_),
    .A2(_05863_),
    .B1(_05880_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _24101_ (.A(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .B(_05828_),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_0 _24102_ (.A1(net3463),
    .A2(_05828_),
    .B1(_05881_),
    .Y(_01153_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_205 ();
 sky130_fd_sc_hd__nand2_1 _24105_ (.A(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .B(_05863_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21ai_0 _24106_ (.A1(_02145_),
    .A2(_05863_),
    .B1(_05884_),
    .Y(_01154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_204 ();
 sky130_fd_sc_hd__nand2_1 _24108_ (.A(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .B(_05863_),
    .Y(_05886_));
 sky130_fd_sc_hd__o21ai_0 _24109_ (.A1(_02297_),
    .A2(_05863_),
    .B1(_05886_),
    .Y(_01155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_203 ();
 sky130_fd_sc_hd__nand2_1 _24111_ (.A(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .B(_05863_),
    .Y(_05888_));
 sky130_fd_sc_hd__o21ai_0 _24112_ (.A1(_02414_),
    .A2(_05863_),
    .B1(_05888_),
    .Y(_01156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_202 ();
 sky130_fd_sc_hd__nand2_1 _24114_ (.A(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .B(_05863_),
    .Y(_05890_));
 sky130_fd_sc_hd__o21ai_0 _24115_ (.A1(_02535_),
    .A2(_05863_),
    .B1(_05890_),
    .Y(_01157_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_200 ();
 sky130_fd_sc_hd__nand2_1 _24118_ (.A(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .B(_05863_),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_0 _24119_ (.A1(_02628_),
    .A2(_05863_),
    .B1(_05893_),
    .Y(_01158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_199 ();
 sky130_fd_sc_hd__nand2_1 _24121_ (.A(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .B(_05863_),
    .Y(_05895_));
 sky130_fd_sc_hd__o21ai_0 _24122_ (.A1(net3453),
    .A2(_05863_),
    .B1(_05895_),
    .Y(_01159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_198 ();
 sky130_fd_sc_hd__nand2_1 _24124_ (.A(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .B(_05863_),
    .Y(_05897_));
 sky130_fd_sc_hd__o21ai_0 _24125_ (.A1(_02837_),
    .A2(_05863_),
    .B1(_05897_),
    .Y(_01160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_197 ();
 sky130_fd_sc_hd__nand2_1 _24127_ (.A(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .B(_05863_),
    .Y(_05899_));
 sky130_fd_sc_hd__o21ai_0 _24128_ (.A1(_02963_),
    .A2(_05863_),
    .B1(_05899_),
    .Y(_01161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_196 ();
 sky130_fd_sc_hd__nand2_1 _24130_ (.A(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .B(_05863_),
    .Y(_05901_));
 sky130_fd_sc_hd__o21ai_0 _24131_ (.A1(net3447),
    .A2(_05863_),
    .B1(_05901_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_4 _24132_ (.A(_05147_),
    .B(_05841_),
    .Y(_05902_));
 sky130_fd_sc_hd__nand2_1 _24133_ (.A(net3446),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_1 _24134_ (.A(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .B(_05863_),
    .Y(_05904_));
 sky130_fd_sc_hd__nand2_1 _24135_ (.A(_05903_),
    .B(_05904_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _24136_ (.A(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .B(_05828_),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_0 _24137_ (.A1(net3459),
    .A2(_05828_),
    .B1(_05905_),
    .Y(_01164_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_195 ();
 sky130_fd_sc_hd__nand2_1 _24139_ (.A(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .B(_05863_),
    .Y(_05907_));
 sky130_fd_sc_hd__o21ai_0 _24140_ (.A1(net3425),
    .A2(_05863_),
    .B1(_05907_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _24141_ (.A(net3416),
    .B(_05902_),
    .Y(_05908_));
 sky130_fd_sc_hd__nand2_1 _24142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .B(_05863_),
    .Y(_05909_));
 sky130_fd_sc_hd__nand2_1 _24143_ (.A(_05908_),
    .B(_05909_),
    .Y(_01166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_194 ();
 sky130_fd_sc_hd__nand2_1 _24145_ (.A(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .B(_05863_),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_0 _24146_ (.A1(net3433),
    .A2(_05863_),
    .B1(_05911_),
    .Y(_01167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_193 ();
 sky130_fd_sc_hd__nand2_1 _24148_ (.A(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .B(_05863_),
    .Y(_05913_));
 sky130_fd_sc_hd__o21ai_0 _24149_ (.A1(net3413),
    .A2(_05863_),
    .B1(_05913_),
    .Y(_01168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_192 ();
 sky130_fd_sc_hd__mux2_1 _24151_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A1(net3412),
    .S(_05902_),
    .X(_01169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_191 ();
 sky130_fd_sc_hd__nand2_1 _24153_ (.A(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .B(_05863_),
    .Y(_05916_));
 sky130_fd_sc_hd__o21ai_0 _24154_ (.A1(net3411),
    .A2(_05863_),
    .B1(_05916_),
    .Y(_01170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_190 ();
 sky130_fd_sc_hd__nand2_1 _24156_ (.A(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .B(_05863_),
    .Y(_05918_));
 sky130_fd_sc_hd__o21ai_0 _24157_ (.A1(net3410),
    .A2(_05863_),
    .B1(_05918_),
    .Y(_01171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_189 ();
 sky130_fd_sc_hd__nand2_1 _24159_ (.A(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .B(_05863_),
    .Y(_05920_));
 sky130_fd_sc_hd__o21ai_0 _24160_ (.A1(net3409),
    .A2(_05863_),
    .B1(_05920_),
    .Y(_01172_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_188 ();
 sky130_fd_sc_hd__nand2_1 _24162_ (.A(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .B(_05863_),
    .Y(_05922_));
 sky130_fd_sc_hd__o21ai_0 _24163_ (.A1(net3408),
    .A2(_05863_),
    .B1(_05922_),
    .Y(_01173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_187 ();
 sky130_fd_sc_hd__nand2_1 _24165_ (.A(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .B(_05863_),
    .Y(_05924_));
 sky130_fd_sc_hd__o21ai_0 _24166_ (.A1(net3407),
    .A2(_05863_),
    .B1(_05924_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _24167_ (.A(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .B(_05828_),
    .Y(_05925_));
 sky130_fd_sc_hd__o21ai_0 _24168_ (.A1(_04483_),
    .A2(_05828_),
    .B1(_05925_),
    .Y(_01175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_186 ();
 sky130_fd_sc_hd__nand2_1 _24170_ (.A(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .B(_05863_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_0 _24171_ (.A1(net3406),
    .A2(_05863_),
    .B1(_05927_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _24172_ (.A(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .B(_05902_),
    .Y(_05928_));
 sky130_fd_sc_hd__a31oi_1 _24173_ (.A1(net3405),
    .A2(net3457),
    .A3(_05902_),
    .B1(_05928_),
    .Y(_01177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_185 ();
 sky130_fd_sc_hd__mux2_1 _24175_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A1(net3404),
    .S(_05902_),
    .X(_01178_));
 sky130_fd_sc_hd__nor2_1 _24176_ (.A(net3464),
    .B(_05863_),
    .Y(_05930_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_184 ();
 sky130_fd_sc_hd__a22o_1 _24178_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A2(_05863_),
    .B1(_05930_),
    .B2(net3403),
    .X(_01179_));
 sky130_fd_sc_hd__nand2_8 _24179_ (.A(_05165_),
    .B(_05810_),
    .Y(_05932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_181 ();
 sky130_fd_sc_hd__nand2_1 _24183_ (.A(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .B(_05932_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_0 _24184_ (.A1(_05011_),
    .A2(_05932_),
    .B1(_05936_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _24185_ (.A(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .B(_05932_),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_0 _24186_ (.A1(net3456),
    .A2(_05932_),
    .B1(_05937_),
    .Y(_01181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_180 ();
 sky130_fd_sc_hd__nand2_1 _24188_ (.A(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .B(_05932_),
    .Y(_05939_));
 sky130_fd_sc_hd__o21ai_0 _24189_ (.A1(_05059_),
    .A2(_05932_),
    .B1(_05939_),
    .Y(_01182_));
 sky130_fd_sc_hd__nand2_1 _24190_ (.A(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .B(_05932_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21ai_0 _24191_ (.A1(net3463),
    .A2(_05932_),
    .B1(_05940_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _24192_ (.A(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .B(_05932_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_0 _24193_ (.A1(net3459),
    .A2(_05932_),
    .B1(_05941_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _24194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .B(_05932_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21ai_0 _24195_ (.A1(net3451),
    .A2(_05932_),
    .B1(_05942_),
    .Y(_01185_));
 sky130_fd_sc_hd__nand2_1 _24196_ (.A(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .B(_05828_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_0 _24197_ (.A1(net3444),
    .A2(_05828_),
    .B1(_05943_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _24198_ (.A(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .B(_05932_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21ai_0 _24199_ (.A1(net3444),
    .A2(_05932_),
    .B1(_05944_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _24200_ (.A(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .B(_05932_),
    .Y(_05945_));
 sky130_fd_sc_hd__o21ai_0 _24201_ (.A1(_04964_),
    .A2(_05932_),
    .B1(_05945_),
    .Y(_01188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_179 ();
 sky130_fd_sc_hd__nand2_1 _24203_ (.A(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .B(_05932_),
    .Y(_05947_));
 sky130_fd_sc_hd__o21ai_0 _24204_ (.A1(_02145_),
    .A2(_05932_),
    .B1(_05947_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _24205_ (.A(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .B(_05932_),
    .Y(_05948_));
 sky130_fd_sc_hd__o21ai_0 _24206_ (.A1(_02297_),
    .A2(_05932_),
    .B1(_05948_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _24207_ (.A(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .B(_05932_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21ai_0 _24208_ (.A1(_02414_),
    .A2(_05932_),
    .B1(_05949_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .B(_05932_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21ai_0 _24210_ (.A1(_02535_),
    .A2(_05932_),
    .B1(_05950_),
    .Y(_01192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_178 ();
 sky130_fd_sc_hd__nand2_1 _24212_ (.A(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .B(_05932_),
    .Y(_05952_));
 sky130_fd_sc_hd__o21ai_0 _24213_ (.A1(_02628_),
    .A2(_05932_),
    .B1(_05952_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _24214_ (.A(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .B(_05932_),
    .Y(_05953_));
 sky130_fd_sc_hd__o21ai_0 _24215_ (.A1(net3453),
    .A2(_05932_),
    .B1(_05953_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _24216_ (.A(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .B(_05932_),
    .Y(_05954_));
 sky130_fd_sc_hd__o21ai_0 _24217_ (.A1(_02837_),
    .A2(_05932_),
    .B1(_05954_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _24218_ (.A(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .B(_05932_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_0 _24219_ (.A1(_02963_),
    .A2(_05932_),
    .B1(_05955_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _24220_ (.A(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .B(_05828_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_0 _24221_ (.A1(_04964_),
    .A2(_05828_),
    .B1(_05956_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_1 _24222_ (.A(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .B(_05932_),
    .Y(_05957_));
 sky130_fd_sc_hd__o21ai_0 _24223_ (.A1(net3447),
    .A2(_05932_),
    .B1(_05957_),
    .Y(_01198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_177 ();
 sky130_fd_sc_hd__nor2_4 _24225_ (.A(_05191_),
    .B(_05841_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2_1 _24226_ (.A(net3446),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__nand2_1 _24227_ (.A(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .B(_05932_),
    .Y(_05961_));
 sky130_fd_sc_hd__nand2_1 _24228_ (.A(_05960_),
    .B(_05961_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _24229_ (.A(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .B(_05932_),
    .Y(_05962_));
 sky130_fd_sc_hd__o21ai_0 _24230_ (.A1(net3425),
    .A2(_05932_),
    .B1(_05962_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _24231_ (.A(net3416),
    .B(_05959_),
    .Y(_05963_));
 sky130_fd_sc_hd__nand2_1 _24232_ (.A(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .B(_05932_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2_1 _24233_ (.A(_05963_),
    .B(_05964_),
    .Y(_01201_));
 sky130_fd_sc_hd__nand2_1 _24234_ (.A(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .B(_05932_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21ai_0 _24235_ (.A1(net3433),
    .A2(_05932_),
    .B1(_05965_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _24236_ (.A(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .B(_05932_),
    .Y(_05966_));
 sky130_fd_sc_hd__o21ai_0 _24237_ (.A1(net3413),
    .A2(_05932_),
    .B1(_05966_),
    .Y(_01203_));
 sky130_fd_sc_hd__mux2_1 _24238_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .A1(net3412),
    .S(_05959_),
    .X(_01204_));
 sky130_fd_sc_hd__nand2_1 _24239_ (.A(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .B(_05932_),
    .Y(_05967_));
 sky130_fd_sc_hd__o21ai_0 _24240_ (.A1(net3411),
    .A2(_05932_),
    .B1(_05967_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _24241_ (.A(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .B(_05932_),
    .Y(_05968_));
 sky130_fd_sc_hd__o21ai_0 _24242_ (.A1(net3410),
    .A2(_05932_),
    .B1(_05968_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _24243_ (.A(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .B(_05932_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21ai_0 _24244_ (.A1(net3409),
    .A2(_05932_),
    .B1(_05969_),
    .Y(_01207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_176 ();
 sky130_fd_sc_hd__nand2_1 _24246_ (.A(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .B(_05828_),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_0 _24247_ (.A1(_02145_),
    .A2(_05828_),
    .B1(_05971_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_1 _24248_ (.A(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .B(_05932_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_0 _24249_ (.A1(net3408),
    .A2(_05932_),
    .B1(_05972_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _24250_ (.A(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .B(_05932_),
    .Y(_05973_));
 sky130_fd_sc_hd__o21ai_0 _24251_ (.A1(net3407),
    .A2(_05932_),
    .B1(_05973_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _24252_ (.A(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .B(_05932_),
    .Y(_05974_));
 sky130_fd_sc_hd__o21ai_0 _24253_ (.A1(net3406),
    .A2(_05932_),
    .B1(_05974_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _24254_ (.A(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .B(_05959_),
    .Y(_05975_));
 sky130_fd_sc_hd__a31oi_1 _24255_ (.A1(net3405),
    .A2(net3457),
    .A3(_05959_),
    .B1(_05975_),
    .Y(_01212_));
 sky130_fd_sc_hd__mux2_1 _24256_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .A1(net3404),
    .S(_05959_),
    .X(_01213_));
 sky130_fd_sc_hd__nor2_1 _24257_ (.A(net3464),
    .B(_05932_),
    .Y(_05976_));
 sky130_fd_sc_hd__a22o_1 _24258_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A2(_05932_),
    .B1(_05976_),
    .B2(net3403),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_8 _24259_ (.A(_02151_),
    .B(_05810_),
    .Y(_05977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_173 ();
 sky130_fd_sc_hd__nand2_1 _24263_ (.A(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .B(_05977_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_0 _24264_ (.A1(_05011_),
    .A2(_05977_),
    .B1(_05981_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand2_1 _24265_ (.A(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .B(_05977_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_0 _24266_ (.A1(net3456),
    .A2(_05977_),
    .B1(_05982_),
    .Y(_01216_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_172 ();
 sky130_fd_sc_hd__nand2_1 _24268_ (.A(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .B(_05977_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21ai_0 _24269_ (.A1(_05059_),
    .A2(_05977_),
    .B1(_05984_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_1 _24270_ (.A(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .B(_05977_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_0 _24271_ (.A1(net3463),
    .A2(_05977_),
    .B1(_05985_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand2_1 _24272_ (.A(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .B(_05828_),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_0 _24273_ (.A1(_02297_),
    .A2(_05828_),
    .B1(_05986_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _24274_ (.A(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .B(_05977_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_0 _24275_ (.A1(net3459),
    .A2(_05977_),
    .B1(_05987_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_1 _24276_ (.A(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .B(_05977_),
    .Y(_05988_));
 sky130_fd_sc_hd__o21ai_0 _24277_ (.A1(net3451),
    .A2(_05977_),
    .B1(_05988_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _24278_ (.A(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .B(_05977_),
    .Y(_05989_));
 sky130_fd_sc_hd__o21ai_0 _24279_ (.A1(net3444),
    .A2(_05977_),
    .B1(_05989_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _24280_ (.A(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .B(_05977_),
    .Y(_05990_));
 sky130_fd_sc_hd__o21ai_0 _24281_ (.A1(_04964_),
    .A2(_05977_),
    .B1(_05990_),
    .Y(_01223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_171 ();
 sky130_fd_sc_hd__nand2_1 _24283_ (.A(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .B(_05977_),
    .Y(_05992_));
 sky130_fd_sc_hd__o21ai_0 _24284_ (.A1(_02145_),
    .A2(_05977_),
    .B1(_05992_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2_1 _24285_ (.A(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .B(_05977_),
    .Y(_05993_));
 sky130_fd_sc_hd__o21ai_0 _24286_ (.A1(_02297_),
    .A2(_05977_),
    .B1(_05993_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _24287_ (.A(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .B(_05977_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21ai_0 _24288_ (.A1(_02414_),
    .A2(_05977_),
    .B1(_05994_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand2_1 _24289_ (.A(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .B(_05977_),
    .Y(_05995_));
 sky130_fd_sc_hd__o21ai_0 _24290_ (.A1(_02535_),
    .A2(_05977_),
    .B1(_05995_),
    .Y(_01227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_170 ();
 sky130_fd_sc_hd__nand2_1 _24292_ (.A(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .B(_05977_),
    .Y(_05997_));
 sky130_fd_sc_hd__o21ai_0 _24293_ (.A1(_02628_),
    .A2(_05977_),
    .B1(_05997_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _24294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .B(_05977_),
    .Y(_05998_));
 sky130_fd_sc_hd__o21ai_0 _24295_ (.A1(net3453),
    .A2(_05977_),
    .B1(_05998_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _24296_ (.A(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .B(_05828_),
    .Y(_05999_));
 sky130_fd_sc_hd__o21ai_0 _24297_ (.A1(_02414_),
    .A2(_05828_),
    .B1(_05999_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _24298_ (.A(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .B(_05977_),
    .Y(_06000_));
 sky130_fd_sc_hd__o21ai_0 _24299_ (.A1(_02837_),
    .A2(_05977_),
    .B1(_06000_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _24300_ (.A(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .B(_05977_),
    .Y(_06001_));
 sky130_fd_sc_hd__o21ai_0 _24301_ (.A1(_02963_),
    .A2(_05977_),
    .B1(_06001_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _24302_ (.A(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .B(_05977_),
    .Y(_06002_));
 sky130_fd_sc_hd__o21ai_0 _24303_ (.A1(net3447),
    .A2(_05977_),
    .B1(_06002_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_4 _24304_ (.A(_03094_),
    .B(_05841_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _24305_ (.A(net3446),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2_1 _24306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .B(_05977_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2_1 _24307_ (.A(_06004_),
    .B(_06005_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand2_1 _24308_ (.A(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .B(_05977_),
    .Y(_06006_));
 sky130_fd_sc_hd__o21ai_0 _24309_ (.A1(net3425),
    .A2(_05977_),
    .B1(_06006_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_1 _24310_ (.A(net3416),
    .B(_06003_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand2_1 _24311_ (.A(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .B(_05977_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _24312_ (.A(_06007_),
    .B(_06008_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _24313_ (.A(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .B(_05977_),
    .Y(_06009_));
 sky130_fd_sc_hd__o21ai_0 _24314_ (.A1(net3433),
    .A2(_05977_),
    .B1(_06009_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _24315_ (.A(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .B(_05977_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21ai_0 _24316_ (.A1(net3413),
    .A2(_05977_),
    .B1(_06010_),
    .Y(_01238_));
 sky130_fd_sc_hd__mux2_1 _24317_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .A1(net3412),
    .S(_06003_),
    .X(_01239_));
 sky130_fd_sc_hd__nand2_1 _24318_ (.A(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .B(_05977_),
    .Y(_06011_));
 sky130_fd_sc_hd__o21ai_0 _24319_ (.A1(net3411),
    .A2(_05977_),
    .B1(_06011_),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .B(_05828_),
    .Y(_06012_));
 sky130_fd_sc_hd__o21ai_0 _24321_ (.A1(_02535_),
    .A2(_05828_),
    .B1(_06012_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _24322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .B(_05977_),
    .Y(_06013_));
 sky130_fd_sc_hd__o21ai_0 _24323_ (.A1(net3410),
    .A2(_05977_),
    .B1(_06013_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_1 _24324_ (.A(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .B(_05977_),
    .Y(_06014_));
 sky130_fd_sc_hd__o21ai_0 _24325_ (.A1(net3409),
    .A2(_05977_),
    .B1(_06014_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _24326_ (.A(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .B(_05977_),
    .Y(_06015_));
 sky130_fd_sc_hd__o21ai_0 _24327_ (.A1(net3408),
    .A2(_05977_),
    .B1(_06015_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2_1 _24328_ (.A(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .B(_05977_),
    .Y(_06016_));
 sky130_fd_sc_hd__o21ai_0 _24329_ (.A1(net3407),
    .A2(_05977_),
    .B1(_06016_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _24330_ (.A(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .B(_05977_),
    .Y(_06017_));
 sky130_fd_sc_hd__o21ai_0 _24331_ (.A1(net3406),
    .A2(_05977_),
    .B1(_06017_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _24332_ (.A(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .B(_06003_),
    .Y(_06018_));
 sky130_fd_sc_hd__a31oi_1 _24333_ (.A1(net3405),
    .A2(net3457),
    .A3(_06003_),
    .B1(_06018_),
    .Y(_01247_));
 sky130_fd_sc_hd__mux2_1 _24334_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .A1(net3404),
    .S(_06003_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _24335_ (.A(net3464),
    .B(_05977_),
    .Y(_06019_));
 sky130_fd_sc_hd__a22o_1 _24336_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .A2(_05977_),
    .B1(_06019_),
    .B2(net3403),
    .X(_01249_));
 sky130_fd_sc_hd__and3b_4 _24337_ (.A_N(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .X(_06020_));
 sky130_fd_sc_hd__nand2_8 _24338_ (.A(_05015_),
    .B(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_167 ();
 sky130_fd_sc_hd__nand2_1 _24342_ (.A(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .B(_06021_),
    .Y(_06025_));
 sky130_fd_sc_hd__o21ai_0 _24343_ (.A1(_05011_),
    .A2(_06021_),
    .B1(_06025_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _24344_ (.A(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .B(_06021_),
    .Y(_06026_));
 sky130_fd_sc_hd__o21ai_0 _24345_ (.A1(_05039_),
    .A2(_06021_),
    .B1(_06026_),
    .Y(_01251_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_166 ();
 sky130_fd_sc_hd__nand2_1 _24347_ (.A(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .B(_05828_),
    .Y(_06028_));
 sky130_fd_sc_hd__o21ai_0 _24348_ (.A1(_02628_),
    .A2(_05828_),
    .B1(_06028_),
    .Y(_01252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_165 ();
 sky130_fd_sc_hd__nand2_1 _24350_ (.A(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .B(_06021_),
    .Y(_06030_));
 sky130_fd_sc_hd__o21ai_0 _24351_ (.A1(_05059_),
    .A2(_06021_),
    .B1(_06030_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _24352_ (.A(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .B(_06021_),
    .Y(_06031_));
 sky130_fd_sc_hd__o21ai_0 _24353_ (.A1(net3463),
    .A2(_06021_),
    .B1(_06031_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _24354_ (.A(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .B(_06021_),
    .Y(_06032_));
 sky130_fd_sc_hd__o21ai_0 _24355_ (.A1(net3459),
    .A2(_06021_),
    .B1(_06032_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _24356_ (.A(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .B(_06021_),
    .Y(_06033_));
 sky130_fd_sc_hd__o21ai_0 _24357_ (.A1(net3451),
    .A2(_06021_),
    .B1(_06033_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _24358_ (.A(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .B(_06021_),
    .Y(_06034_));
 sky130_fd_sc_hd__o21ai_0 _24359_ (.A1(net3444),
    .A2(_06021_),
    .B1(_06034_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _24360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .B(_06021_),
    .Y(_06035_));
 sky130_fd_sc_hd__o21ai_0 _24361_ (.A1(_04964_),
    .A2(_06021_),
    .B1(_06035_),
    .Y(_01258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_164 ();
 sky130_fd_sc_hd__nand2_1 _24363_ (.A(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .B(_06021_),
    .Y(_06037_));
 sky130_fd_sc_hd__o21ai_0 _24364_ (.A1(_02145_),
    .A2(_06021_),
    .B1(_06037_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _24365_ (.A(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .B(_06021_),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_0 _24366_ (.A1(_02297_),
    .A2(_06021_),
    .B1(_06038_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _24367_ (.A(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .B(_06021_),
    .Y(_06039_));
 sky130_fd_sc_hd__o21ai_0 _24368_ (.A1(_02414_),
    .A2(_06021_),
    .B1(_06039_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2_1 _24369_ (.A(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .B(_06021_),
    .Y(_06040_));
 sky130_fd_sc_hd__o21ai_0 _24370_ (.A1(net3460),
    .A2(_06021_),
    .B1(_06040_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _24371_ (.A(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .B(_05828_),
    .Y(_06041_));
 sky130_fd_sc_hd__o21ai_0 _24372_ (.A1(net3453),
    .A2(_05828_),
    .B1(_06041_),
    .Y(_01263_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_163 ();
 sky130_fd_sc_hd__nand2_1 _24374_ (.A(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .B(_06021_),
    .Y(_06043_));
 sky130_fd_sc_hd__o21ai_0 _24375_ (.A1(_02628_),
    .A2(_06021_),
    .B1(_06043_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _24376_ (.A(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .B(_06021_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21ai_0 _24377_ (.A1(net3453),
    .A2(_06021_),
    .B1(_06044_),
    .Y(_01265_));
 sky130_fd_sc_hd__nand2_1 _24378_ (.A(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .B(_06021_),
    .Y(_06045_));
 sky130_fd_sc_hd__o21ai_0 _24379_ (.A1(_02837_),
    .A2(_06021_),
    .B1(_06045_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _24380_ (.A(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .B(_06021_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21ai_0 _24381_ (.A1(_02963_),
    .A2(_06021_),
    .B1(_06046_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _24382_ (.A(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .B(_06021_),
    .Y(_06047_));
 sky130_fd_sc_hd__o21ai_0 _24383_ (.A1(net3447),
    .A2(_06021_),
    .B1(_06047_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand3b_1 _24384_ (.A_N(net3827),
    .B(net3945),
    .C(net3946),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_4 _24385_ (.A(_05100_),
    .B(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _24386_ (.A(net3446),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_1 _24387_ (.A(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .B(_06021_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _24388_ (.A(_06050_),
    .B(_06051_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_1 _24389_ (.A(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .B(_06021_),
    .Y(_06052_));
 sky130_fd_sc_hd__o21ai_0 _24390_ (.A1(net3425),
    .A2(_06021_),
    .B1(_06052_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _24391_ (.A(net3416),
    .B(_06049_),
    .Y(_06053_));
 sky130_fd_sc_hd__nand2_1 _24392_ (.A(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .B(_06021_),
    .Y(_06054_));
 sky130_fd_sc_hd__nand2_1 _24393_ (.A(_06053_),
    .B(_06054_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _24394_ (.A(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .B(_06021_),
    .Y(_06055_));
 sky130_fd_sc_hd__o21ai_0 _24395_ (.A1(net3433),
    .A2(_06021_),
    .B1(_06055_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _24396_ (.A(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .B(_06021_),
    .Y(_06056_));
 sky130_fd_sc_hd__o21ai_0 _24397_ (.A1(net3413),
    .A2(_06021_),
    .B1(_06056_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _24398_ (.A(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .B(_05828_),
    .Y(_06057_));
 sky130_fd_sc_hd__o21ai_0 _24399_ (.A1(_02837_),
    .A2(_05828_),
    .B1(_06057_),
    .Y(_01274_));
 sky130_fd_sc_hd__mux2_1 _24400_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(net3412),
    .S(_06049_),
    .X(_01275_));
 sky130_fd_sc_hd__nand2_1 _24401_ (.A(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .B(_06021_),
    .Y(_06058_));
 sky130_fd_sc_hd__o21ai_0 _24402_ (.A1(net3411),
    .A2(_06021_),
    .B1(_06058_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _24403_ (.A(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .B(_06021_),
    .Y(_06059_));
 sky130_fd_sc_hd__o21ai_0 _24404_ (.A1(net3410),
    .A2(_06021_),
    .B1(_06059_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _24405_ (.A(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .B(_06021_),
    .Y(_06060_));
 sky130_fd_sc_hd__o21ai_0 _24406_ (.A1(net3409),
    .A2(_06021_),
    .B1(_06060_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _24407_ (.A(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .B(_06021_),
    .Y(_06061_));
 sky130_fd_sc_hd__o21ai_0 _24408_ (.A1(net3408),
    .A2(_06021_),
    .B1(_06061_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2_1 _24409_ (.A(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .B(_06021_),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_0 _24410_ (.A1(net3407),
    .A2(_06021_),
    .B1(_06062_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _24411_ (.A(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .B(_06021_),
    .Y(_06063_));
 sky130_fd_sc_hd__o21ai_0 _24412_ (.A1(net3406),
    .A2(_06021_),
    .B1(_06063_),
    .Y(_01281_));
 sky130_fd_sc_hd__nor2_1 _24413_ (.A(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .B(_06049_),
    .Y(_06064_));
 sky130_fd_sc_hd__a31oi_1 _24414_ (.A1(net3405),
    .A2(net3457),
    .A3(_06049_),
    .B1(_06064_),
    .Y(_01282_));
 sky130_fd_sc_hd__mux2_1 _24415_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(net3404),
    .S(_06049_),
    .X(_01283_));
 sky130_fd_sc_hd__nor2_1 _24416_ (.A(_04920_),
    .B(_06021_),
    .Y(_06065_));
 sky130_fd_sc_hd__a22o_1 _24417_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A2(_06021_),
    .B1(_06065_),
    .B2(net3403),
    .X(_01284_));
 sky130_fd_sc_hd__nand2_1 _24418_ (.A(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .B(_05828_),
    .Y(_06066_));
 sky130_fd_sc_hd__o21ai_0 _24419_ (.A1(_02963_),
    .A2(_05828_),
    .B1(_06066_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_8 _24420_ (.A(_05122_),
    .B(_06020_),
    .Y(_06067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_160 ();
 sky130_fd_sc_hd__nand2_1 _24424_ (.A(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .B(_06067_),
    .Y(_06071_));
 sky130_fd_sc_hd__o21ai_0 _24425_ (.A1(_05011_),
    .A2(_06067_),
    .B1(_06071_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _24426_ (.A(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .B(_06067_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21ai_0 _24427_ (.A1(_05039_),
    .A2(_06067_),
    .B1(_06072_),
    .Y(_01287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_159 ();
 sky130_fd_sc_hd__nand2_1 _24429_ (.A(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .B(_06067_),
    .Y(_06074_));
 sky130_fd_sc_hd__o21ai_0 _24430_ (.A1(_05059_),
    .A2(_06067_),
    .B1(_06074_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _24431_ (.A(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .B(_06067_),
    .Y(_06075_));
 sky130_fd_sc_hd__o21ai_0 _24432_ (.A1(net3463),
    .A2(_06067_),
    .B1(_06075_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _24433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .B(_06067_),
    .Y(_06076_));
 sky130_fd_sc_hd__o21ai_0 _24434_ (.A1(net3459),
    .A2(_06067_),
    .B1(_06076_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _24435_ (.A(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .B(_06067_),
    .Y(_06077_));
 sky130_fd_sc_hd__o21ai_0 _24436_ (.A1(net3451),
    .A2(_06067_),
    .B1(_06077_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand2_1 _24437_ (.A(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .B(_06067_),
    .Y(_06078_));
 sky130_fd_sc_hd__o21ai_0 _24438_ (.A1(net3444),
    .A2(_06067_),
    .B1(_06078_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _24439_ (.A(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .B(_06067_),
    .Y(_06079_));
 sky130_fd_sc_hd__o21ai_0 _24440_ (.A1(_04964_),
    .A2(_06067_),
    .B1(_06079_),
    .Y(_01293_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_158 ();
 sky130_fd_sc_hd__nand2_1 _24442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .B(_06067_),
    .Y(_06081_));
 sky130_fd_sc_hd__o21ai_0 _24443_ (.A1(_02145_),
    .A2(_06067_),
    .B1(_06081_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _24444_ (.A(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .B(_06067_),
    .Y(_06082_));
 sky130_fd_sc_hd__o21ai_0 _24445_ (.A1(_02297_),
    .A2(_06067_),
    .B1(_06082_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _24446_ (.A(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .B(_05828_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_0 _24447_ (.A1(net3447),
    .A2(_05828_),
    .B1(_06083_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _24448_ (.A(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .B(_06067_),
    .Y(_06084_));
 sky130_fd_sc_hd__o21ai_0 _24449_ (.A1(_02414_),
    .A2(_06067_),
    .B1(_06084_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _24450_ (.A(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .B(_06067_),
    .Y(_06085_));
 sky130_fd_sc_hd__o21ai_0 _24451_ (.A1(net3460),
    .A2(_06067_),
    .B1(_06085_),
    .Y(_01298_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_157 ();
 sky130_fd_sc_hd__nand2_1 _24453_ (.A(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .B(_06067_),
    .Y(_06087_));
 sky130_fd_sc_hd__o21ai_0 _24454_ (.A1(_02628_),
    .A2(_06067_),
    .B1(_06087_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _24455_ (.A(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .B(_06067_),
    .Y(_06088_));
 sky130_fd_sc_hd__o21ai_0 _24456_ (.A1(net3453),
    .A2(_06067_),
    .B1(_06088_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _24457_ (.A(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .B(_06067_),
    .Y(_06089_));
 sky130_fd_sc_hd__o21ai_0 _24458_ (.A1(_02837_),
    .A2(_06067_),
    .B1(_06089_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _24459_ (.A(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .B(_06067_),
    .Y(_06090_));
 sky130_fd_sc_hd__o21ai_0 _24460_ (.A1(_02963_),
    .A2(_06067_),
    .B1(_06090_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _24461_ (.A(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .B(_06067_),
    .Y(_06091_));
 sky130_fd_sc_hd__o21ai_0 _24462_ (.A1(net3447),
    .A2(_06067_),
    .B1(_06091_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_4 _24463_ (.A(_05147_),
    .B(_06048_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _24464_ (.A(net3446),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__nand2_1 _24465_ (.A(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .B(_06067_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_1 _24466_ (.A(_06093_),
    .B(_06094_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _24467_ (.A(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .B(_06067_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21ai_0 _24468_ (.A1(net3425),
    .A2(_06067_),
    .B1(_06095_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _24469_ (.A(net3416),
    .B(_06092_),
    .Y(_06096_));
 sky130_fd_sc_hd__nand2_1 _24470_ (.A(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .B(_06067_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _24471_ (.A(_06096_),
    .B(_06097_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_4 _24472_ (.A(_04978_),
    .B(_05191_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _24473_ (.A(net3446),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand2_1 _24474_ (.A(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .B(_05828_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_1 _24475_ (.A(_06099_),
    .B(_06100_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .B(_06067_),
    .Y(_06101_));
 sky130_fd_sc_hd__o21ai_0 _24477_ (.A1(net3433),
    .A2(_06067_),
    .B1(_06101_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_1 _24478_ (.A(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .B(_06067_),
    .Y(_06102_));
 sky130_fd_sc_hd__o21ai_0 _24479_ (.A1(net3413),
    .A2(_06067_),
    .B1(_06102_),
    .Y(_01309_));
 sky130_fd_sc_hd__mux2_1 _24480_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A1(net3412),
    .S(_06092_),
    .X(_01310_));
 sky130_fd_sc_hd__nand2_1 _24481_ (.A(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .B(_06067_),
    .Y(_06103_));
 sky130_fd_sc_hd__o21ai_0 _24482_ (.A1(net3411),
    .A2(_06067_),
    .B1(_06103_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _24483_ (.A(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .B(_06067_),
    .Y(_06104_));
 sky130_fd_sc_hd__o21ai_0 _24484_ (.A1(net3410),
    .A2(_06067_),
    .B1(_06104_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand2_1 _24485_ (.A(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .B(_06067_),
    .Y(_06105_));
 sky130_fd_sc_hd__o21ai_0 _24486_ (.A1(net3409),
    .A2(_06067_),
    .B1(_06105_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _24487_ (.A(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .B(_06067_),
    .Y(_06106_));
 sky130_fd_sc_hd__o21ai_0 _24488_ (.A1(net3408),
    .A2(_06067_),
    .B1(_06106_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _24489_ (.A(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .B(_06067_),
    .Y(_06107_));
 sky130_fd_sc_hd__o21ai_0 _24490_ (.A1(net3407),
    .A2(_06067_),
    .B1(_06107_),
    .Y(_01315_));
 sky130_fd_sc_hd__nand2_1 _24491_ (.A(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .B(_06067_),
    .Y(_06108_));
 sky130_fd_sc_hd__o21ai_0 _24492_ (.A1(net3406),
    .A2(_06067_),
    .B1(_06108_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor2_1 _24493_ (.A(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .B(_06092_),
    .Y(_06109_));
 sky130_fd_sc_hd__a31oi_1 _24494_ (.A1(net3405),
    .A2(net3457),
    .A3(_06092_),
    .B1(_06109_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _24495_ (.A(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .B(_05828_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21ai_0 _24496_ (.A1(net3425),
    .A2(_05828_),
    .B1(_06110_),
    .Y(_01318_));
 sky130_fd_sc_hd__mux2_1 _24497_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A1(net3404),
    .S(_06092_),
    .X(_01319_));
 sky130_fd_sc_hd__nor2_1 _24498_ (.A(_04920_),
    .B(_06067_),
    .Y(_06111_));
 sky130_fd_sc_hd__a22o_1 _24499_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(_06067_),
    .B1(_06111_),
    .B2(net3403),
    .X(_01320_));
 sky130_fd_sc_hd__nand2_8 _24500_ (.A(_05165_),
    .B(_06020_),
    .Y(_06112_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_154 ();
 sky130_fd_sc_hd__nand2_1 _24504_ (.A(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .B(_06112_),
    .Y(_06116_));
 sky130_fd_sc_hd__o21ai_0 _24505_ (.A1(_05011_),
    .A2(_06112_),
    .B1(_06116_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_1 _24506_ (.A(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .B(_06112_),
    .Y(_06117_));
 sky130_fd_sc_hd__o21ai_0 _24507_ (.A1(_05039_),
    .A2(_06112_),
    .B1(_06117_),
    .Y(_01322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_153 ();
 sky130_fd_sc_hd__nand2_1 _24509_ (.A(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .B(_06112_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_0 _24510_ (.A1(_05059_),
    .A2(_06112_),
    .B1(_06119_),
    .Y(_01323_));
 sky130_fd_sc_hd__nand2_1 _24511_ (.A(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .B(_06112_),
    .Y(_06120_));
 sky130_fd_sc_hd__o21ai_0 _24512_ (.A1(net3463),
    .A2(_06112_),
    .B1(_06120_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_1 _24513_ (.A(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .B(_06112_),
    .Y(_06121_));
 sky130_fd_sc_hd__o21ai_0 _24514_ (.A1(net3459),
    .A2(_06112_),
    .B1(_06121_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _24515_ (.A(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .B(_06112_),
    .Y(_06122_));
 sky130_fd_sc_hd__o21ai_0 _24516_ (.A1(net3451),
    .A2(_06112_),
    .B1(_06122_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _24517_ (.A(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .B(_06112_),
    .Y(_06123_));
 sky130_fd_sc_hd__o21ai_0 _24518_ (.A1(net3444),
    .A2(_06112_),
    .B1(_06123_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_1 _24519_ (.A(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .B(_06112_),
    .Y(_06124_));
 sky130_fd_sc_hd__o21ai_0 _24520_ (.A1(_04964_),
    .A2(_06112_),
    .B1(_06124_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _24521_ (.A(net3416),
    .B(_06098_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _24522_ (.A(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .B(_05828_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_1 _24523_ (.A(_06125_),
    .B(_06126_),
    .Y(_01329_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_152 ();
 sky130_fd_sc_hd__nand2_1 _24525_ (.A(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .B(_06112_),
    .Y(_06128_));
 sky130_fd_sc_hd__o21ai_0 _24526_ (.A1(_02145_),
    .A2(_06112_),
    .B1(_06128_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _24527_ (.A(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .B(_06112_),
    .Y(_06129_));
 sky130_fd_sc_hd__o21ai_0 _24528_ (.A1(_02297_),
    .A2(_06112_),
    .B1(_06129_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _24529_ (.A(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .B(_06112_),
    .Y(_06130_));
 sky130_fd_sc_hd__o21ai_0 _24530_ (.A1(_02414_),
    .A2(_06112_),
    .B1(_06130_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _24531_ (.A(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .B(_06112_),
    .Y(_06131_));
 sky130_fd_sc_hd__o21ai_0 _24532_ (.A1(net3460),
    .A2(_06112_),
    .B1(_06131_),
    .Y(_01333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_151 ();
 sky130_fd_sc_hd__nand2_1 _24534_ (.A(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .B(_06112_),
    .Y(_06133_));
 sky130_fd_sc_hd__o21ai_0 _24535_ (.A1(_02628_),
    .A2(_06112_),
    .B1(_06133_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_1 _24536_ (.A(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .B(_06112_),
    .Y(_06134_));
 sky130_fd_sc_hd__o21ai_0 _24537_ (.A1(net3453),
    .A2(_06112_),
    .B1(_06134_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _24538_ (.A(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .B(_06112_),
    .Y(_06135_));
 sky130_fd_sc_hd__o21ai_0 _24539_ (.A1(_02837_),
    .A2(_06112_),
    .B1(_06135_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _24540_ (.A(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .B(_06112_),
    .Y(_06136_));
 sky130_fd_sc_hd__o21ai_0 _24541_ (.A1(_02963_),
    .A2(_06112_),
    .B1(_06136_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _24542_ (.A(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .B(_06112_),
    .Y(_06137_));
 sky130_fd_sc_hd__o21ai_0 _24543_ (.A1(net3447),
    .A2(_06112_),
    .B1(_06137_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_4 _24544_ (.A(_05191_),
    .B(_06048_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2_1 _24545_ (.A(net3446),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__nand2_1 _24546_ (.A(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .B(_06112_),
    .Y(_06140_));
 sky130_fd_sc_hd__nand2_1 _24547_ (.A(_06139_),
    .B(_06140_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2_1 _24548_ (.A(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .B(_05828_),
    .Y(_06141_));
 sky130_fd_sc_hd__o21ai_0 _24549_ (.A1(net3433),
    .A2(_05828_),
    .B1(_06141_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _24550_ (.A(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .B(_06112_),
    .Y(_06142_));
 sky130_fd_sc_hd__o21ai_0 _24551_ (.A1(net3425),
    .A2(_06112_),
    .B1(_06142_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_1 _24552_ (.A(net3416),
    .B(_06138_),
    .Y(_06143_));
 sky130_fd_sc_hd__nand2_1 _24553_ (.A(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .B(_06112_),
    .Y(_06144_));
 sky130_fd_sc_hd__nand2_1 _24554_ (.A(_06143_),
    .B(_06144_),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _24555_ (.A(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .B(_06112_),
    .Y(_06145_));
 sky130_fd_sc_hd__o21ai_0 _24556_ (.A1(net3433),
    .A2(_06112_),
    .B1(_06145_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _24557_ (.A(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .B(_06112_),
    .Y(_06146_));
 sky130_fd_sc_hd__o21ai_0 _24558_ (.A1(net3413),
    .A2(_06112_),
    .B1(_06146_),
    .Y(_01344_));
 sky130_fd_sc_hd__mux2_1 _24559_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A1(net3412),
    .S(_06138_),
    .X(_01345_));
 sky130_fd_sc_hd__nand2_1 _24560_ (.A(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .B(_06112_),
    .Y(_06147_));
 sky130_fd_sc_hd__o21ai_0 _24561_ (.A1(net3411),
    .A2(_06112_),
    .B1(_06147_),
    .Y(_01346_));
 sky130_fd_sc_hd__nand2_1 _24562_ (.A(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .B(_06112_),
    .Y(_06148_));
 sky130_fd_sc_hd__o21ai_0 _24563_ (.A1(net3410),
    .A2(_06112_),
    .B1(_06148_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _24564_ (.A(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .B(_06112_),
    .Y(_06149_));
 sky130_fd_sc_hd__o21ai_0 _24565_ (.A1(net3409),
    .A2(_06112_),
    .B1(_06149_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _24566_ (.A(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .B(_06112_),
    .Y(_06150_));
 sky130_fd_sc_hd__o21ai_0 _24567_ (.A1(net3408),
    .A2(_06112_),
    .B1(_06150_),
    .Y(_01349_));
 sky130_fd_sc_hd__nand2_1 _24568_ (.A(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .B(_06112_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21ai_0 _24569_ (.A1(net3407),
    .A2(_06112_),
    .B1(_06151_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _24570_ (.A(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .B(_05828_),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_0 _24571_ (.A1(net3413),
    .A2(_05828_),
    .B1(_06152_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_1 _24572_ (.A(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .B(_06112_),
    .Y(_06153_));
 sky130_fd_sc_hd__o21ai_0 _24573_ (.A1(net3406),
    .A2(_06112_),
    .B1(_06153_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _24574_ (.A(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .B(_06138_),
    .Y(_06154_));
 sky130_fd_sc_hd__a31oi_1 _24575_ (.A1(net3405),
    .A2(net3457),
    .A3(_06138_),
    .B1(_06154_),
    .Y(_01353_));
 sky130_fd_sc_hd__mux2_1 _24576_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A1(net3404),
    .S(_06138_),
    .X(_01354_));
 sky130_fd_sc_hd__nor2_1 _24577_ (.A(_04920_),
    .B(_06112_),
    .Y(_06155_));
 sky130_fd_sc_hd__a22o_1 _24578_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A2(_06112_),
    .B1(_06155_),
    .B2(net3403),
    .X(_01355_));
 sky130_fd_sc_hd__nand2_8 _24579_ (.A(_02151_),
    .B(_06020_),
    .Y(_06156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_148 ();
 sky130_fd_sc_hd__nand2_1 _24583_ (.A(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .B(_06156_),
    .Y(_06160_));
 sky130_fd_sc_hd__o21ai_0 _24584_ (.A1(_05011_),
    .A2(_06156_),
    .B1(_06160_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _24585_ (.A(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .B(_06156_),
    .Y(_06161_));
 sky130_fd_sc_hd__o21ai_0 _24586_ (.A1(_05039_),
    .A2(_06156_),
    .B1(_06161_),
    .Y(_01357_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_147 ();
 sky130_fd_sc_hd__nand2_1 _24588_ (.A(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .B(_06156_),
    .Y(_06163_));
 sky130_fd_sc_hd__o21ai_0 _24589_ (.A1(_05059_),
    .A2(_06156_),
    .B1(_06163_),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_1 _24590_ (.A(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .B(_06156_),
    .Y(_06164_));
 sky130_fd_sc_hd__o21ai_0 _24591_ (.A1(net3463),
    .A2(_06156_),
    .B1(_06164_),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_1 _24592_ (.A(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .B(_06156_),
    .Y(_06165_));
 sky130_fd_sc_hd__o21ai_0 _24593_ (.A1(net3459),
    .A2(_06156_),
    .B1(_06165_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _24594_ (.A(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .B(_06156_),
    .Y(_06166_));
 sky130_fd_sc_hd__o21ai_0 _24595_ (.A1(net3451),
    .A2(_06156_),
    .B1(_06166_),
    .Y(_01361_));
 sky130_fd_sc_hd__mux2_1 _24596_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A1(net3412),
    .S(_06098_),
    .X(_01362_));
 sky130_fd_sc_hd__nand2_1 _24597_ (.A(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .B(_06156_),
    .Y(_06167_));
 sky130_fd_sc_hd__o21ai_0 _24598_ (.A1(net3444),
    .A2(_06156_),
    .B1(_06167_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _24599_ (.A(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .B(_06156_),
    .Y(_06168_));
 sky130_fd_sc_hd__o21ai_0 _24600_ (.A1(_04964_),
    .A2(_06156_),
    .B1(_06168_),
    .Y(_01364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_146 ();
 sky130_fd_sc_hd__nand2_1 _24602_ (.A(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .B(_06156_),
    .Y(_06170_));
 sky130_fd_sc_hd__o21ai_0 _24603_ (.A1(_02145_),
    .A2(_06156_),
    .B1(_06170_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _24604_ (.A(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .B(_06156_),
    .Y(_06171_));
 sky130_fd_sc_hd__o21ai_0 _24605_ (.A1(_02297_),
    .A2(_06156_),
    .B1(_06171_),
    .Y(_01366_));
 sky130_fd_sc_hd__nand2_1 _24606_ (.A(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .B(_06156_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21ai_0 _24607_ (.A1(_02414_),
    .A2(_06156_),
    .B1(_06172_),
    .Y(_01367_));
 sky130_fd_sc_hd__nand2_1 _24608_ (.A(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .B(_06156_),
    .Y(_06173_));
 sky130_fd_sc_hd__o21ai_0 _24609_ (.A1(net3460),
    .A2(_06156_),
    .B1(_06173_),
    .Y(_01368_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_145 ();
 sky130_fd_sc_hd__nand2_1 _24611_ (.A(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .B(_06156_),
    .Y(_06175_));
 sky130_fd_sc_hd__o21ai_0 _24612_ (.A1(_02628_),
    .A2(_06156_),
    .B1(_06175_),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2_1 _24613_ (.A(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .B(_06156_),
    .Y(_06176_));
 sky130_fd_sc_hd__o21ai_0 _24614_ (.A1(net3453),
    .A2(_06156_),
    .B1(_06176_),
    .Y(_01370_));
 sky130_fd_sc_hd__nand2_1 _24615_ (.A(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .B(_06156_),
    .Y(_06177_));
 sky130_fd_sc_hd__o21ai_0 _24616_ (.A1(_02837_),
    .A2(_06156_),
    .B1(_06177_),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2_1 _24617_ (.A(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .B(_06156_),
    .Y(_06178_));
 sky130_fd_sc_hd__o21ai_0 _24618_ (.A1(_02963_),
    .A2(_06156_),
    .B1(_06178_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _24619_ (.A(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .B(_05828_),
    .Y(_06179_));
 sky130_fd_sc_hd__o21ai_0 _24620_ (.A1(net3411),
    .A2(_05828_),
    .B1(_06179_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _24621_ (.A(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .B(_06156_),
    .Y(_06180_));
 sky130_fd_sc_hd__o21ai_0 _24622_ (.A1(net3447),
    .A2(_06156_),
    .B1(_06180_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_4 _24623_ (.A(_03094_),
    .B(_06048_),
    .Y(_06181_));
 sky130_fd_sc_hd__nand2_1 _24624_ (.A(net3446),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _24625_ (.A(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .B(_06156_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_1 _24626_ (.A(_06182_),
    .B(_06183_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _24627_ (.A(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .B(_06156_),
    .Y(_06184_));
 sky130_fd_sc_hd__o21ai_0 _24628_ (.A1(net3425),
    .A2(_06156_),
    .B1(_06184_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _24629_ (.A(net3416),
    .B(_06181_),
    .Y(_06185_));
 sky130_fd_sc_hd__nand2_1 _24630_ (.A(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .B(_06156_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _24631_ (.A(_06185_),
    .B(_06186_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _24632_ (.A(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .B(_06156_),
    .Y(_06187_));
 sky130_fd_sc_hd__o21ai_0 _24633_ (.A1(net3433),
    .A2(_06156_),
    .B1(_06187_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _24634_ (.A(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .B(_06156_),
    .Y(_06188_));
 sky130_fd_sc_hd__o21ai_0 _24635_ (.A1(net3413),
    .A2(_06156_),
    .B1(_06188_),
    .Y(_01379_));
 sky130_fd_sc_hd__mux2_1 _24636_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .A1(net3412),
    .S(_06181_),
    .X(_01380_));
 sky130_fd_sc_hd__nand2_1 _24637_ (.A(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .B(_06156_),
    .Y(_06189_));
 sky130_fd_sc_hd__o21ai_0 _24638_ (.A1(net3411),
    .A2(_06156_),
    .B1(_06189_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _24639_ (.A(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .B(_06156_),
    .Y(_06190_));
 sky130_fd_sc_hd__o21ai_0 _24640_ (.A1(net3410),
    .A2(_06156_),
    .B1(_06190_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _24641_ (.A(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .B(_06156_),
    .Y(_06191_));
 sky130_fd_sc_hd__o21ai_0 _24642_ (.A1(net3409),
    .A2(_06156_),
    .B1(_06191_),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2_1 _24643_ (.A(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .B(_05828_),
    .Y(_06192_));
 sky130_fd_sc_hd__o21ai_0 _24644_ (.A1(net3410),
    .A2(_05828_),
    .B1(_06192_),
    .Y(_01384_));
 sky130_fd_sc_hd__nand2_1 _24645_ (.A(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .B(_06156_),
    .Y(_06193_));
 sky130_fd_sc_hd__o21ai_0 _24646_ (.A1(net3408),
    .A2(_06156_),
    .B1(_06193_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _24647_ (.A(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .B(_06156_),
    .Y(_06194_));
 sky130_fd_sc_hd__o21ai_0 _24648_ (.A1(net3407),
    .A2(_06156_),
    .B1(_06194_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _24649_ (.A(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .B(_06156_),
    .Y(_06195_));
 sky130_fd_sc_hd__o21ai_0 _24650_ (.A1(net3406),
    .A2(_06156_),
    .B1(_06195_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _24651_ (.A(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .B(_06181_),
    .Y(_06196_));
 sky130_fd_sc_hd__a31oi_1 _24652_ (.A1(net3405),
    .A2(net3457),
    .A3(_06181_),
    .B1(_06196_),
    .Y(_01388_));
 sky130_fd_sc_hd__mux2_1 _24653_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .A1(net3404),
    .S(_06181_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_1 _24654_ (.A(_04920_),
    .B(_06156_),
    .Y(_06197_));
 sky130_fd_sc_hd__a22o_1 _24655_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .A2(_06156_),
    .B1(_06197_),
    .B2(net3403),
    .X(_01390_));
 sky130_fd_sc_hd__nand2_8 _24656_ (.A(_02147_),
    .B(_05015_),
    .Y(_06198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__nand2_1 _24660_ (.A(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .B(_06198_),
    .Y(_06202_));
 sky130_fd_sc_hd__o21ai_0 _24661_ (.A1(_05011_),
    .A2(_06198_),
    .B1(_06202_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _24662_ (.A(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .B(_06198_),
    .Y(_06203_));
 sky130_fd_sc_hd__o21ai_0 _24663_ (.A1(_05039_),
    .A2(_06198_),
    .B1(_06203_),
    .Y(_01392_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__nand2_1 _24665_ (.A(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .B(_06198_),
    .Y(_06205_));
 sky130_fd_sc_hd__o21ai_0 _24666_ (.A1(_05059_),
    .A2(_06198_),
    .B1(_06205_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2_1 _24667_ (.A(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .B(_06198_),
    .Y(_06206_));
 sky130_fd_sc_hd__o21ai_0 _24668_ (.A1(net3463),
    .A2(_06198_),
    .B1(_06206_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _24669_ (.A(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .B(_05828_),
    .Y(_06207_));
 sky130_fd_sc_hd__o21ai_0 _24670_ (.A1(net3409),
    .A2(_05828_),
    .B1(_06207_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _24671_ (.A(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .B(_06198_),
    .Y(_06208_));
 sky130_fd_sc_hd__o21ai_0 _24672_ (.A1(net3459),
    .A2(_06198_),
    .B1(_06208_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _24673_ (.A(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .B(_06198_),
    .Y(_06209_));
 sky130_fd_sc_hd__o21ai_0 _24674_ (.A1(net3451),
    .A2(_06198_),
    .B1(_06209_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _24675_ (.A(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .B(_06198_),
    .Y(_06210_));
 sky130_fd_sc_hd__o21ai_0 _24676_ (.A1(net3444),
    .A2(_06198_),
    .B1(_06210_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _24677_ (.A(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .B(_06198_),
    .Y(_06211_));
 sky130_fd_sc_hd__o21ai_0 _24678_ (.A1(_04964_),
    .A2(_06198_),
    .B1(_06211_),
    .Y(_01399_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__nand2_1 _24680_ (.A(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .B(_06198_),
    .Y(_06213_));
 sky130_fd_sc_hd__o21ai_0 _24681_ (.A1(_02145_),
    .A2(_06198_),
    .B1(_06213_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_1 _24682_ (.A(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .B(_06198_),
    .Y(_06214_));
 sky130_fd_sc_hd__o21ai_0 _24683_ (.A1(_02297_),
    .A2(_06198_),
    .B1(_06214_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand2_1 _24684_ (.A(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .B(_06198_),
    .Y(_06215_));
 sky130_fd_sc_hd__o21ai_0 _24685_ (.A1(_02414_),
    .A2(_06198_),
    .B1(_06215_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_1 _24686_ (.A(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .B(_06198_),
    .Y(_06216_));
 sky130_fd_sc_hd__o21ai_0 _24687_ (.A1(net3460),
    .A2(_06198_),
    .B1(_06216_),
    .Y(_01403_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__nand2_1 _24689_ (.A(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .B(_06198_),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_0 _24690_ (.A1(_02628_),
    .A2(_06198_),
    .B1(_06218_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _24691_ (.A(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .B(_06198_),
    .Y(_06219_));
 sky130_fd_sc_hd__o21ai_0 _24692_ (.A1(net3453),
    .A2(_06198_),
    .B1(_06219_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand2_1 _24693_ (.A(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .B(_05828_),
    .Y(_06220_));
 sky130_fd_sc_hd__o21ai_0 _24694_ (.A1(net3408),
    .A2(_05828_),
    .B1(_06220_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _24695_ (.A(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .B(_06198_),
    .Y(_06221_));
 sky130_fd_sc_hd__o21ai_0 _24696_ (.A1(_02837_),
    .A2(_06198_),
    .B1(_06221_),
    .Y(_01407_));
 sky130_fd_sc_hd__nand2_1 _24697_ (.A(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .B(_06198_),
    .Y(_06222_));
 sky130_fd_sc_hd__o21ai_0 _24698_ (.A1(_02963_),
    .A2(_06198_),
    .B1(_06222_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _24699_ (.A(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .B(_06198_),
    .Y(_06223_));
 sky130_fd_sc_hd__o21ai_0 _24700_ (.A1(net3447),
    .A2(_06198_),
    .B1(_06223_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_4 _24701_ (.A(_03093_),
    .B(_05100_),
    .Y(_06224_));
 sky130_fd_sc_hd__nand2_1 _24702_ (.A(net3446),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__nand2_1 _24703_ (.A(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .B(_06198_),
    .Y(_06226_));
 sky130_fd_sc_hd__nand2_1 _24704_ (.A(_06225_),
    .B(_06226_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_1 _24705_ (.A(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .B(_06198_),
    .Y(_06227_));
 sky130_fd_sc_hd__o21ai_0 _24706_ (.A1(net3425),
    .A2(_06198_),
    .B1(_06227_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _24707_ (.A(net3416),
    .B(_06224_),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_1 _24708_ (.A(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .B(_06198_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2_1 _24709_ (.A(_06228_),
    .B(_06229_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _24710_ (.A(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .B(_06198_),
    .Y(_06230_));
 sky130_fd_sc_hd__o21ai_0 _24711_ (.A1(net3433),
    .A2(_06198_),
    .B1(_06230_),
    .Y(_01413_));
 sky130_fd_sc_hd__nand2_1 _24712_ (.A(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .B(_06198_),
    .Y(_06231_));
 sky130_fd_sc_hd__o21ai_0 _24713_ (.A1(net3413),
    .A2(_06198_),
    .B1(_06231_),
    .Y(_01414_));
 sky130_fd_sc_hd__mux2_1 _24714_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A1(net3412),
    .S(_06224_),
    .X(_01415_));
 sky130_fd_sc_hd__nand2_1 _24715_ (.A(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .B(_06198_),
    .Y(_06232_));
 sky130_fd_sc_hd__o21ai_0 _24716_ (.A1(net3411),
    .A2(_06198_),
    .B1(_06232_),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2_1 _24717_ (.A(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .B(_05828_),
    .Y(_06233_));
 sky130_fd_sc_hd__o21ai_0 _24718_ (.A1(net3407),
    .A2(_05828_),
    .B1(_06233_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _24719_ (.A(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .B(_06198_),
    .Y(_06234_));
 sky130_fd_sc_hd__o21ai_0 _24720_ (.A1(net3410),
    .A2(_06198_),
    .B1(_06234_),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2_1 _24721_ (.A(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .B(_06198_),
    .Y(_06235_));
 sky130_fd_sc_hd__o21ai_0 _24722_ (.A1(net3409),
    .A2(_06198_),
    .B1(_06235_),
    .Y(_01419_));
 sky130_fd_sc_hd__nand2_1 _24723_ (.A(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .B(_06198_),
    .Y(_06236_));
 sky130_fd_sc_hd__o21ai_0 _24724_ (.A1(net3408),
    .A2(_06198_),
    .B1(_06236_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _24725_ (.A(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .B(_06198_),
    .Y(_06237_));
 sky130_fd_sc_hd__o21ai_0 _24726_ (.A1(net3407),
    .A2(_06198_),
    .B1(_06237_),
    .Y(_01421_));
 sky130_fd_sc_hd__nand2_1 _24727_ (.A(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .B(_06198_),
    .Y(_06238_));
 sky130_fd_sc_hd__o21ai_0 _24728_ (.A1(net3406),
    .A2(_06198_),
    .B1(_06238_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _24729_ (.A(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .B(_06224_),
    .Y(_06239_));
 sky130_fd_sc_hd__a31oi_1 _24730_ (.A1(net3405),
    .A2(net3457),
    .A3(_06224_),
    .B1(_06239_),
    .Y(_01423_));
 sky130_fd_sc_hd__mux2_1 _24731_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A1(net3404),
    .S(_06224_),
    .X(_01424_));
 sky130_fd_sc_hd__nor2_1 _24732_ (.A(_04920_),
    .B(_06198_),
    .Y(_06240_));
 sky130_fd_sc_hd__a22o_1 _24733_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A2(_06198_),
    .B1(_06240_),
    .B2(net3403),
    .X(_01425_));
 sky130_fd_sc_hd__nand2_8 _24734_ (.A(_02147_),
    .B(_05122_),
    .Y(_06241_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_136 ();
 sky130_fd_sc_hd__nand2_1 _24738_ (.A(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .B(_06241_),
    .Y(_06245_));
 sky130_fd_sc_hd__o21ai_0 _24739_ (.A1(_05011_),
    .A2(_06241_),
    .B1(_06245_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _24740_ (.A(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .B(_06241_),
    .Y(_06246_));
 sky130_fd_sc_hd__o21ai_0 _24741_ (.A1(_05039_),
    .A2(_06241_),
    .B1(_06246_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _24742_ (.A(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .B(_05828_),
    .Y(_06247_));
 sky130_fd_sc_hd__o21ai_0 _24743_ (.A1(net3406),
    .A2(_05828_),
    .B1(_06247_),
    .Y(_01428_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__nand2_1 _24745_ (.A(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .B(_06241_),
    .Y(_06249_));
 sky130_fd_sc_hd__o21ai_0 _24746_ (.A1(_05059_),
    .A2(_06241_),
    .B1(_06249_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _24747_ (.A(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .B(_06241_),
    .Y(_06250_));
 sky130_fd_sc_hd__o21ai_0 _24748_ (.A1(net3463),
    .A2(_06241_),
    .B1(_06250_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _24749_ (.A(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .B(_06241_),
    .Y(_06251_));
 sky130_fd_sc_hd__o21ai_0 _24750_ (.A1(net3459),
    .A2(_06241_),
    .B1(_06251_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _24751_ (.A(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .B(_06241_),
    .Y(_06252_));
 sky130_fd_sc_hd__o21ai_0 _24752_ (.A1(net3451),
    .A2(_06241_),
    .B1(_06252_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _24753_ (.A(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .B(_06241_),
    .Y(_06253_));
 sky130_fd_sc_hd__o21ai_0 _24754_ (.A1(net3444),
    .A2(_06241_),
    .B1(_06253_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _24755_ (.A(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .B(_06241_),
    .Y(_06254_));
 sky130_fd_sc_hd__o21ai_0 _24756_ (.A1(_04964_),
    .A2(_06241_),
    .B1(_06254_),
    .Y(_01434_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__nand2_1 _24758_ (.A(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .B(_06241_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21ai_0 _24759_ (.A1(_02145_),
    .A2(_06241_),
    .B1(_06256_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _24760_ (.A(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .B(_06241_),
    .Y(_06257_));
 sky130_fd_sc_hd__o21ai_0 _24761_ (.A1(_02297_),
    .A2(_06241_),
    .B1(_06257_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _24762_ (.A(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .B(_06241_),
    .Y(_06258_));
 sky130_fd_sc_hd__o21ai_0 _24763_ (.A1(_02414_),
    .A2(_06241_),
    .B1(_06258_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _24764_ (.A(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .B(_06241_),
    .Y(_06259_));
 sky130_fd_sc_hd__o21ai_0 _24765_ (.A1(net3460),
    .A2(_06241_),
    .B1(_06259_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _24766_ (.A(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .B(_06098_),
    .Y(_06260_));
 sky130_fd_sc_hd__a31oi_1 _24767_ (.A1(net3405),
    .A2(net3457),
    .A3(_06098_),
    .B1(_06260_),
    .Y(_01439_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_133 ();
 sky130_fd_sc_hd__nand2_1 _24769_ (.A(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .B(_06241_),
    .Y(_06262_));
 sky130_fd_sc_hd__o21ai_0 _24770_ (.A1(_02628_),
    .A2(_06241_),
    .B1(_06262_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_1 _24771_ (.A(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .B(_06241_),
    .Y(_06263_));
 sky130_fd_sc_hd__o21ai_0 _24772_ (.A1(net3453),
    .A2(_06241_),
    .B1(_06263_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _24773_ (.A(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .B(_06241_),
    .Y(_06264_));
 sky130_fd_sc_hd__o21ai_0 _24774_ (.A1(_02837_),
    .A2(_06241_),
    .B1(_06264_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _24775_ (.A(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .B(_06241_),
    .Y(_06265_));
 sky130_fd_sc_hd__o21ai_0 _24776_ (.A1(_02963_),
    .A2(_06241_),
    .B1(_06265_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _24777_ (.A(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .B(_06241_),
    .Y(_06266_));
 sky130_fd_sc_hd__o21ai_0 _24778_ (.A1(net3447),
    .A2(_06241_),
    .B1(_06266_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_4 _24779_ (.A(_03093_),
    .B(_05147_),
    .Y(_06267_));
 sky130_fd_sc_hd__nand2_1 _24780_ (.A(net3446),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _24781_ (.A(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .B(_06241_),
    .Y(_06269_));
 sky130_fd_sc_hd__nand2_1 _24782_ (.A(_06268_),
    .B(_06269_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _24783_ (.A(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .B(_06241_),
    .Y(_06270_));
 sky130_fd_sc_hd__o21ai_0 _24784_ (.A1(net3425),
    .A2(_06241_),
    .B1(_06270_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _24785_ (.A(net3416),
    .B(_06267_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_1 _24786_ (.A(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .B(_06241_),
    .Y(_06272_));
 sky130_fd_sc_hd__nand2_1 _24787_ (.A(_06271_),
    .B(_06272_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _24788_ (.A(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .B(_06241_),
    .Y(_06273_));
 sky130_fd_sc_hd__o21ai_0 _24789_ (.A1(net3433),
    .A2(_06241_),
    .B1(_06273_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _24790_ (.A(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .B(_06241_),
    .Y(_06274_));
 sky130_fd_sc_hd__o21ai_0 _24791_ (.A1(net3413),
    .A2(_06241_),
    .B1(_06274_),
    .Y(_01449_));
 sky130_fd_sc_hd__mux2_1 _24792_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A1(net3404),
    .S(_06098_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _24793_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A1(net3412),
    .S(_06267_),
    .X(_01451_));
 sky130_fd_sc_hd__nand2_1 _24794_ (.A(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .B(_06241_),
    .Y(_06275_));
 sky130_fd_sc_hd__o21ai_0 _24795_ (.A1(net3411),
    .A2(_06241_),
    .B1(_06275_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_1 _24796_ (.A(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .B(_06241_),
    .Y(_06276_));
 sky130_fd_sc_hd__o21ai_0 _24797_ (.A1(net3410),
    .A2(_06241_),
    .B1(_06276_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _24798_ (.A(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .B(_06241_),
    .Y(_06277_));
 sky130_fd_sc_hd__o21ai_0 _24799_ (.A1(net3409),
    .A2(_06241_),
    .B1(_06277_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _24800_ (.A(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .B(_06241_),
    .Y(_06278_));
 sky130_fd_sc_hd__o21ai_0 _24801_ (.A1(net3408),
    .A2(_06241_),
    .B1(_06278_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _24802_ (.A(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .B(_06241_),
    .Y(_06279_));
 sky130_fd_sc_hd__o21ai_0 _24803_ (.A1(net3407),
    .A2(_06241_),
    .B1(_06279_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _24804_ (.A(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .B(_06241_),
    .Y(_06280_));
 sky130_fd_sc_hd__o21ai_0 _24805_ (.A1(net3406),
    .A2(_06241_),
    .B1(_06280_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _24806_ (.A(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .B(_06267_),
    .Y(_06281_));
 sky130_fd_sc_hd__a31oi_1 _24807_ (.A1(net3405),
    .A2(net3457),
    .A3(_06267_),
    .B1(_06281_),
    .Y(_01458_));
 sky130_fd_sc_hd__mux2_1 _24808_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A1(net3404),
    .S(_06267_),
    .X(_01459_));
 sky130_fd_sc_hd__nor2_1 _24809_ (.A(_04920_),
    .B(_06241_),
    .Y(_06282_));
 sky130_fd_sc_hd__a22o_1 _24810_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(_06241_),
    .B1(_06282_),
    .B2(net3403),
    .X(_01460_));
 sky130_fd_sc_hd__nor2_1 _24811_ (.A(_04920_),
    .B(_05828_),
    .Y(_06283_));
 sky130_fd_sc_hd__a22o_1 _24812_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(_05828_),
    .B1(_06283_),
    .B2(net3403),
    .X(_01461_));
 sky130_fd_sc_hd__nand2_8 _24813_ (.A(_02147_),
    .B(_05165_),
    .Y(_06284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_130 ();
 sky130_fd_sc_hd__nand2_1 _24817_ (.A(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .B(_06284_),
    .Y(_06288_));
 sky130_fd_sc_hd__o21ai_0 _24818_ (.A1(_05011_),
    .A2(_06284_),
    .B1(_06288_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _24819_ (.A(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .B(_06284_),
    .Y(_06289_));
 sky130_fd_sc_hd__o21ai_0 _24820_ (.A1(_05039_),
    .A2(_06284_),
    .B1(_06289_),
    .Y(_01463_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_129 ();
 sky130_fd_sc_hd__nand2_1 _24822_ (.A(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .B(_06284_),
    .Y(_06291_));
 sky130_fd_sc_hd__o21ai_0 _24823_ (.A1(_05059_),
    .A2(_06284_),
    .B1(_06291_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _24824_ (.A(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .B(_06284_),
    .Y(_06292_));
 sky130_fd_sc_hd__o21ai_0 _24825_ (.A1(net3463),
    .A2(_06284_),
    .B1(_06292_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _24826_ (.A(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .B(_06284_),
    .Y(_06293_));
 sky130_fd_sc_hd__o21ai_0 _24827_ (.A1(net3459),
    .A2(_06284_),
    .B1(_06293_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _24828_ (.A(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .B(_06284_),
    .Y(_06294_));
 sky130_fd_sc_hd__o21ai_0 _24829_ (.A1(net3451),
    .A2(_06284_),
    .B1(_06294_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _24830_ (.A(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .B(_06284_),
    .Y(_06295_));
 sky130_fd_sc_hd__o21ai_0 _24831_ (.A1(net3444),
    .A2(_06284_),
    .B1(_06295_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _24832_ (.A(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .B(_06284_),
    .Y(_06296_));
 sky130_fd_sc_hd__o21ai_0 _24833_ (.A1(_04964_),
    .A2(_06284_),
    .B1(_06296_),
    .Y(_01469_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_128 ();
 sky130_fd_sc_hd__nand2_1 _24835_ (.A(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .B(_06284_),
    .Y(_06298_));
 sky130_fd_sc_hd__o21ai_0 _24836_ (.A1(_02145_),
    .A2(_06284_),
    .B1(_06298_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _24837_ (.A(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .B(_06284_),
    .Y(_06299_));
 sky130_fd_sc_hd__o21ai_0 _24838_ (.A1(_02297_),
    .A2(_06284_),
    .B1(_06299_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _24839_ (.A(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .B(_03280_),
    .Y(_06300_));
 sky130_fd_sc_hd__o21ai_0 _24840_ (.A1(_03280_),
    .A2(_05011_),
    .B1(_06300_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _24841_ (.A(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .B(_06284_),
    .Y(_06301_));
 sky130_fd_sc_hd__o21ai_0 _24842_ (.A1(_02414_),
    .A2(_06284_),
    .B1(_06301_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _24843_ (.A(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .B(_06284_),
    .Y(_06302_));
 sky130_fd_sc_hd__o21ai_0 _24844_ (.A1(net3460),
    .A2(_06284_),
    .B1(_06302_),
    .Y(_01474_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_127 ();
 sky130_fd_sc_hd__nand2_1 _24846_ (.A(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .B(_06284_),
    .Y(_06304_));
 sky130_fd_sc_hd__o21ai_0 _24847_ (.A1(_02628_),
    .A2(_06284_),
    .B1(_06304_),
    .Y(_01475_));
 sky130_fd_sc_hd__nand2_1 _24848_ (.A(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .B(_06284_),
    .Y(_06305_));
 sky130_fd_sc_hd__o21ai_0 _24849_ (.A1(net3453),
    .A2(_06284_),
    .B1(_06305_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _24850_ (.A(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .B(_06284_),
    .Y(_06306_));
 sky130_fd_sc_hd__o21ai_0 _24851_ (.A1(_02837_),
    .A2(_06284_),
    .B1(_06306_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _24852_ (.A(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .B(_06284_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21ai_0 _24853_ (.A1(_02963_),
    .A2(_06284_),
    .B1(_06307_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _24854_ (.A(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .B(_06284_),
    .Y(_06308_));
 sky130_fd_sc_hd__o21ai_0 _24855_ (.A1(net3447),
    .A2(_06284_),
    .B1(_06308_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_4 _24856_ (.A(_03093_),
    .B(_05191_),
    .Y(_06309_));
 sky130_fd_sc_hd__nand2_1 _24857_ (.A(net3446),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand2_1 _24858_ (.A(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .B(_06284_),
    .Y(_06311_));
 sky130_fd_sc_hd__nand2_1 _24859_ (.A(_06310_),
    .B(_06311_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _24860_ (.A(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .B(_06284_),
    .Y(_06312_));
 sky130_fd_sc_hd__o21ai_0 _24861_ (.A1(net3425),
    .A2(_06284_),
    .B1(_06312_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_1 _24862_ (.A(net3416),
    .B(_06309_),
    .Y(_06313_));
 sky130_fd_sc_hd__nand2_1 _24863_ (.A(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .B(_06284_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand2_1 _24864_ (.A(_06313_),
    .B(_06314_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _24865_ (.A(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .B(_03280_),
    .Y(_06315_));
 sky130_fd_sc_hd__o21ai_0 _24866_ (.A1(_03280_),
    .A2(_05039_),
    .B1(_06315_),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _24867_ (.A(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .B(_06284_),
    .Y(_06316_));
 sky130_fd_sc_hd__o21ai_0 _24868_ (.A1(net3433),
    .A2(_06284_),
    .B1(_06316_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _24869_ (.A(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .B(_06284_),
    .Y(_06317_));
 sky130_fd_sc_hd__o21ai_0 _24870_ (.A1(net3413),
    .A2(_06284_),
    .B1(_06317_),
    .Y(_01485_));
 sky130_fd_sc_hd__mux2_1 _24871_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .A1(net3412),
    .S(_06309_),
    .X(_01486_));
 sky130_fd_sc_hd__nand2_1 _24872_ (.A(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .B(_06284_),
    .Y(_06318_));
 sky130_fd_sc_hd__o21ai_0 _24873_ (.A1(net3411),
    .A2(_06284_),
    .B1(_06318_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _24874_ (.A(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .B(_06284_),
    .Y(_06319_));
 sky130_fd_sc_hd__o21ai_0 _24875_ (.A1(net3410),
    .A2(_06284_),
    .B1(_06319_),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_1 _24876_ (.A(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .B(_06284_),
    .Y(_06320_));
 sky130_fd_sc_hd__o21ai_0 _24877_ (.A1(net3409),
    .A2(_06284_),
    .B1(_06320_),
    .Y(_01489_));
 sky130_fd_sc_hd__nand2_1 _24878_ (.A(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .B(_06284_),
    .Y(_06321_));
 sky130_fd_sc_hd__o21ai_0 _24879_ (.A1(net3408),
    .A2(_06284_),
    .B1(_06321_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _24880_ (.A(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .B(_06284_),
    .Y(_06322_));
 sky130_fd_sc_hd__o21ai_0 _24881_ (.A1(net3407),
    .A2(_06284_),
    .B1(_06322_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _24882_ (.A(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .B(_06284_),
    .Y(_06323_));
 sky130_fd_sc_hd__o21ai_0 _24883_ (.A1(net3406),
    .A2(_06284_),
    .B1(_06323_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _24884_ (.A(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .B(_06309_),
    .Y(_06324_));
 sky130_fd_sc_hd__a31oi_1 _24885_ (.A1(net3405),
    .A2(net3457),
    .A3(_06309_),
    .B1(_06324_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _24886_ (.A(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .B(_03280_),
    .Y(_06325_));
 sky130_fd_sc_hd__o21ai_0 _24887_ (.A1(_03280_),
    .A2(_05059_),
    .B1(_06325_),
    .Y(_01494_));
 sky130_fd_sc_hd__mux2_1 _24888_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .A1(net3404),
    .S(_06309_),
    .X(_01495_));
 sky130_fd_sc_hd__nor2_1 _24889_ (.A(_04920_),
    .B(_06284_),
    .Y(_06326_));
 sky130_fd_sc_hd__a22o_1 _24890_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A2(_06284_),
    .B1(_06326_),
    .B2(net3403),
    .X(_01496_));
 sky130_fd_sc_hd__nand2_1 _24891_ (.A(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .B(_02153_),
    .Y(_06327_));
 sky130_fd_sc_hd__o21ai_0 _24892_ (.A1(_02153_),
    .A2(_05011_),
    .B1(_06327_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_1 _24893_ (.A(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .B(_02153_),
    .Y(_06328_));
 sky130_fd_sc_hd__o21ai_0 _24894_ (.A1(_02153_),
    .A2(_05039_),
    .B1(_06328_),
    .Y(_01498_));
 sky130_fd_sc_hd__nand2_1 _24895_ (.A(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .B(_02153_),
    .Y(_06329_));
 sky130_fd_sc_hd__o21ai_0 _24896_ (.A1(_02153_),
    .A2(_05059_),
    .B1(_06329_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _24897_ (.A(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .B(_02153_),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ai_0 _24898_ (.A1(_02153_),
    .A2(net3463),
    .B1(_06330_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _24899_ (.A(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .B(_02153_),
    .Y(_06331_));
 sky130_fd_sc_hd__o21ai_0 _24900_ (.A1(_02153_),
    .A2(net3459),
    .B1(_06331_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand2_1 _24901_ (.A(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .B(_02153_),
    .Y(_06332_));
 sky130_fd_sc_hd__o21ai_0 _24902_ (.A1(_02153_),
    .A2(net3451),
    .B1(_06332_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _24903_ (.A(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .B(_02153_),
    .Y(_06333_));
 sky130_fd_sc_hd__o21ai_0 _24904_ (.A1(_02153_),
    .A2(net3444),
    .B1(_06333_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _24905_ (.A(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .B(_02153_),
    .Y(_06334_));
 sky130_fd_sc_hd__o21ai_0 _24906_ (.A1(_02153_),
    .A2(_04964_),
    .B1(_06334_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _24907_ (.A(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .B(_03280_),
    .Y(_06335_));
 sky130_fd_sc_hd__o21ai_0 _24908_ (.A1(_03280_),
    .A2(net3463),
    .B1(_06335_),
    .Y(_01505_));
 sky130_fd_sc_hd__or2_4 _24909_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_10974_),
    .X(_06336_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_126 ();
 sky130_fd_sc_hd__nor2_1 _24911_ (.A(net3448),
    .B(_06336_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _24912_ (.A(_10650_),
    .B(_10972_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor3_1 _24913_ (.A(_10540_),
    .B(_06338_),
    .C(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__o21ai_0 _24914_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_10975_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _24915_ (.A(_10495_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__or2_4 _24916_ (.A(_10504_),
    .B(_10514_),
    .X(_06343_));
 sky130_fd_sc_hd__a41o_4 _24917_ (.A1(net3895),
    .A2(_10646_),
    .A3(_12411_),
    .A4(_10791_),
    .B1(_06336_),
    .X(_06344_));
 sky130_fd_sc_hd__o21ai_2 _24918_ (.A1(_06343_),
    .A2(_10784_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _24919_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_06346_));
 sky130_fd_sc_hd__o21ai_0 _24920_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_06345_),
    .B1(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__nand2_1 _24921_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__a21oi_1 _24922_ (.A1(_06342_),
    .A2(_06348_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Y(_06349_));
 sky130_fd_sc_hd__nor4_1 _24923_ (.A(\cs_registers_i.debug_mode_i ),
    .B(\cs_registers_i.dcsr_q[2] ),
    .C(net60),
    .D(_10821_),
    .Y(_06350_));
 sky130_fd_sc_hd__nor3b_4 _24924_ (.A(_10495_),
    .B(_10978_),
    .C_N(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__nor4_1 _24925_ (.A(_12176_),
    .B(_06340_),
    .C(_06349_),
    .D(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__nor2_1 _24926_ (.A(net3448),
    .B(_10979_),
    .Y(_06353_));
 sky130_fd_sc_hd__nand3_1 _24927_ (.A(_10495_),
    .B(_10539_),
    .C(_06336_),
    .Y(_06354_));
 sky130_fd_sc_hd__nor3_1 _24928_ (.A(_10823_),
    .B(_06353_),
    .C(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__nor2_1 _24929_ (.A(_06352_),
    .B(_06355_),
    .Y(_01506_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_123 ();
 sky130_fd_sc_hd__nand3_1 _24933_ (.A(net3742),
    .B(_10823_),
    .C(_06336_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_1 _24934_ (.A(net3742),
    .B(_06339_),
    .Y(_06360_));
 sky130_fd_sc_hd__o21ai_0 _24935_ (.A1(_12169_),
    .A2(_10970_),
    .B1(_06343_),
    .Y(_06361_));
 sky130_fd_sc_hd__nor3_1 _24936_ (.A(_10500_),
    .B(_10784_),
    .C(_10796_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand3_1 _24937_ (.A(_10539_),
    .B(_10823_),
    .C(_06336_),
    .Y(_06363_));
 sky130_fd_sc_hd__a21oi_1 _24938_ (.A1(_10978_),
    .A2(_06363_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_06364_));
 sky130_fd_sc_hd__a311oi_1 _24939_ (.A1(_06344_),
    .A2(_06361_),
    .A3(_06362_),
    .B1(_06364_),
    .C1(_06351_),
    .Y(_06365_));
 sky130_fd_sc_hd__o211ai_1 _24940_ (.A1(net3448),
    .A2(_06359_),
    .B1(_06360_),
    .C1(_06365_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand3_1 _24941_ (.A(_10650_),
    .B(_10972_),
    .C(_06338_),
    .Y(_06366_));
 sky130_fd_sc_hd__nor3_1 _24942_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10538_),
    .C(_10975_),
    .Y(_06367_));
 sky130_fd_sc_hd__a21oi_1 _24943_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_10977_),
    .B1(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__o21ai_0 _24944_ (.A1(_10498_),
    .A2(_10798_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_06369_));
 sky130_fd_sc_hd__o221ai_1 _24945_ (.A1(_10795_),
    .A2(_06345_),
    .B1(_06368_),
    .B2(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C1(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__a21oi_1 _24946_ (.A1(net3742),
    .A2(_06366_),
    .B1(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__nor2b_1 _24947_ (.A(_10798_),
    .B_N(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Y(_06372_));
 sky130_fd_sc_hd__nor3_1 _24948_ (.A(_06351_),
    .B(_06371_),
    .C(_06372_),
    .Y(_01508_));
 sky130_fd_sc_hd__o21ai_0 _24949_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_06336_),
    .B1(_06366_),
    .Y(_06373_));
 sky130_fd_sc_hd__a21oi_1 _24950_ (.A1(_10794_),
    .A2(_06344_),
    .B1(_10500_),
    .Y(_06374_));
 sky130_fd_sc_hd__a21o_1 _24951_ (.A1(_10539_),
    .A2(_06373_),
    .B1(_06374_),
    .X(_01509_));
 sky130_fd_sc_hd__nor3_1 _24952_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\cs_registers_i.dcsr_q[2] ),
    .C(net60),
    .Y(_06375_));
 sky130_fd_sc_hd__o31ai_1 _24953_ (.A1(_10642_),
    .A2(_12167_),
    .A3(_12176_),
    .B1(\cs_registers_i.debug_mode_i ),
    .Y(_06376_));
 sky130_fd_sc_hd__o21ai_0 _24954_ (.A1(_12171_),
    .A2(_06375_),
    .B1(_06376_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21oi_1 _24955_ (.A1(net145),
    .A2(net3573),
    .B1(\cs_registers_i.nmi_mode_i ),
    .Y(_06377_));
 sky130_fd_sc_hd__nor2_1 _24956_ (.A(net3663),
    .B(_06377_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand3b_1 _24957_ (.A_N(net3753),
    .B(_10779_),
    .C(_10924_),
    .Y(_06378_));
 sky130_fd_sc_hd__a31oi_1 _24958_ (.A1(_07883_),
    .A2(_08040_),
    .A3(_05003_),
    .B1(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_1 _24959_ (.A(_02148_),
    .B(_10657_),
    .Y(_06380_));
 sky130_fd_sc_hd__nand3_1 _24960_ (.A(net3673),
    .B(_10924_),
    .C(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _24961_ (.A(\id_stage_i.id_fsm_q ),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__o21ai_0 _24962_ (.A1(_10780_),
    .A2(_06379_),
    .B1(_06382_),
    .Y(_01512_));
 sky130_fd_sc_hd__mux2_1 _24963_ (.A0(net3712),
    .A1(net3575),
    .S(net3631),
    .X(_06383_));
 sky130_fd_sc_hd__nand2_8 _24964_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_10980_),
    .Y(_06384_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_122 ();
 sky130_fd_sc_hd__nand2_1 _24966_ (.A(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .B(_06384_),
    .Y(_06386_));
 sky130_fd_sc_hd__o21ai_0 _24967_ (.A1(_10684_),
    .A2(_06383_),
    .B1(_06386_),
    .Y(_01513_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_121 ();
 sky130_fd_sc_hd__mux2i_1 _24969_ (.A0(net3515),
    .A1(net3701),
    .S(_04421_),
    .Y(_06388_));
 sky130_fd_sc_hd__nand2_1 _24970_ (.A(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .B(_06384_),
    .Y(_06389_));
 sky130_fd_sc_hd__o21ai_0 _24971_ (.A1(_10684_),
    .A2(_06388_),
    .B1(_06389_),
    .Y(_01514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_120 ();
 sky130_fd_sc_hd__nor2_1 _24973_ (.A(_09030_),
    .B(net3631),
    .Y(_06391_));
 sky130_fd_sc_hd__a21oi_1 _24974_ (.A1(net152),
    .A2(net3631),
    .B1(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_1 _24975_ (.A(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .B(_06384_),
    .Y(_06393_));
 sky130_fd_sc_hd__o21ai_0 _24976_ (.A1(_10684_),
    .A2(_06392_),
    .B1(_06393_),
    .Y(_01515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_119 ();
 sky130_fd_sc_hd__nand2_1 _24978_ (.A(_09243_),
    .B(_02990_),
    .Y(_06395_));
 sky130_fd_sc_hd__o21ai_0 _24979_ (.A1(net3514),
    .A2(_04421_),
    .B1(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand2_1 _24980_ (.A(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .B(_06384_),
    .Y(_06397_));
 sky130_fd_sc_hd__o21ai_0 _24981_ (.A1(_10684_),
    .A2(_06396_),
    .B1(_06397_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _24982_ (.A(_09149_),
    .B(net3631),
    .Y(_06398_));
 sky130_fd_sc_hd__a21oi_1 _24983_ (.A1(net154),
    .A2(net3631),
    .B1(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand2_1 _24984_ (.A(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .B(_06384_),
    .Y(_06400_));
 sky130_fd_sc_hd__o21ai_0 _24985_ (.A1(_10684_),
    .A2(_06399_),
    .B1(_06400_),
    .Y(_01517_));
 sky130_fd_sc_hd__mux2i_1 _24986_ (.A0(net3513),
    .A1(net3696),
    .S(_04421_),
    .Y(_06401_));
 sky130_fd_sc_hd__nand2_1 _24987_ (.A(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .B(_06384_),
    .Y(_06402_));
 sky130_fd_sc_hd__o21ai_0 _24988_ (.A1(_10684_),
    .A2(_06401_),
    .B1(_06402_),
    .Y(_01518_));
 sky130_fd_sc_hd__nand2_1 _24989_ (.A(net389),
    .B(_02990_),
    .Y(_06403_));
 sky130_fd_sc_hd__o21ai_0 _24990_ (.A1(net3507),
    .A2(_02990_),
    .B1(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2_1 _24991_ (.A(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .B(_06384_),
    .Y(_06405_));
 sky130_fd_sc_hd__o21ai_0 _24992_ (.A1(_10684_),
    .A2(_06404_),
    .B1(_06405_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _24993_ (.A(_09512_),
    .B(net3631),
    .Y(_06406_));
 sky130_fd_sc_hd__a21oi_1 _24994_ (.A1(net3506),
    .A2(net3631),
    .B1(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__nand2_1 _24995_ (.A(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .B(_06384_),
    .Y(_06408_));
 sky130_fd_sc_hd__o21ai_0 _24996_ (.A1(_10684_),
    .A2(_06407_),
    .B1(_06408_),
    .Y(_01520_));
 sky130_fd_sc_hd__mux2i_1 _24997_ (.A0(net3512),
    .A1(net409),
    .S(_04421_),
    .Y(_06409_));
 sky130_fd_sc_hd__nand2_1 _24998_ (.A(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .B(_06384_),
    .Y(_06410_));
 sky130_fd_sc_hd__o21ai_0 _24999_ (.A1(_10684_),
    .A2(_06409_),
    .B1(_06410_),
    .Y(_01521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_118 ();
 sky130_fd_sc_hd__nor2_1 _25001_ (.A(net3497),
    .B(_02990_),
    .Y(_06412_));
 sky130_fd_sc_hd__a21oi_1 _25002_ (.A1(net3692),
    .A2(_02990_),
    .B1(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_117 ();
 sky130_fd_sc_hd__nand2_1 _25004_ (.A(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .B(_06384_),
    .Y(_06415_));
 sky130_fd_sc_hd__o21ai_0 _25005_ (.A1(_10684_),
    .A2(_06413_),
    .B1(_06415_),
    .Y(_01522_));
 sky130_fd_sc_hd__mux2i_1 _25006_ (.A0(net160),
    .A1(_09564_),
    .S(_04421_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2_1 _25007_ (.A(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .B(_06384_),
    .Y(_06417_));
 sky130_fd_sc_hd__o21ai_0 _25008_ (.A1(_10684_),
    .A2(_06416_),
    .B1(_06417_),
    .Y(_01523_));
 sky130_fd_sc_hd__xnor2_4 _25009_ (.A(net3583),
    .B(net3574),
    .Y(_06418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_115 ();
 sky130_fd_sc_hd__nand2_1 _25012_ (.A(net342),
    .B(_02990_),
    .Y(_06421_));
 sky130_fd_sc_hd__o21ai_0 _25013_ (.A1(net3556),
    .A2(_04421_),
    .B1(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_1 _25014_ (.A(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .B(_06384_),
    .Y(_06423_));
 sky130_fd_sc_hd__o21ai_0 _25015_ (.A1(_10684_),
    .A2(_06422_),
    .B1(_06423_),
    .Y(_01524_));
 sky130_fd_sc_hd__mux2i_1 _25016_ (.A0(net451),
    .A1(net3688),
    .S(_04421_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand2_1 _25017_ (.A(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .B(_06384_),
    .Y(_06425_));
 sky130_fd_sc_hd__o21ai_0 _25018_ (.A1(_10684_),
    .A2(_06424_),
    .B1(_06425_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor2_1 _25019_ (.A(net3496),
    .B(_02990_),
    .Y(_06426_));
 sky130_fd_sc_hd__a21oi_1 _25020_ (.A1(net3691),
    .A2(_02990_),
    .B1(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _25021_ (.A(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .B(_06384_),
    .Y(_06428_));
 sky130_fd_sc_hd__o21ai_0 _25022_ (.A1(_10684_),
    .A2(_06427_),
    .B1(_06428_),
    .Y(_01526_));
 sky130_fd_sc_hd__mux2i_1 _25023_ (.A0(net3686),
    .A1(net3503),
    .S(net3631),
    .Y(_06429_));
 sky130_fd_sc_hd__nand2_1 _25024_ (.A(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .B(_06384_),
    .Y(_06430_));
 sky130_fd_sc_hd__o21ai_0 _25025_ (.A1(_06384_),
    .A2(_06429_),
    .B1(_06430_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _25026_ (.A(net3504),
    .B(_02990_),
    .Y(_06431_));
 sky130_fd_sc_hd__a21oi_1 _25027_ (.A1(net3685),
    .A2(_02990_),
    .B1(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_1 _25028_ (.A(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .B(_06384_),
    .Y(_06433_));
 sky130_fd_sc_hd__o21ai_0 _25029_ (.A1(_10684_),
    .A2(_06432_),
    .B1(_06433_),
    .Y(_01528_));
 sky130_fd_sc_hd__mux2i_1 _25030_ (.A0(_10010_),
    .A1(net274),
    .S(net3631),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_1 _25031_ (.A(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .B(_06384_),
    .Y(_06435_));
 sky130_fd_sc_hd__o21ai_0 _25032_ (.A1(_06384_),
    .A2(_06434_),
    .B1(_06435_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _25033_ (.A(_10062_),
    .B(net3631),
    .Y(_06436_));
 sky130_fd_sc_hd__a21oi_1 _25034_ (.A1(net3495),
    .A2(net3631),
    .B1(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand2_1 _25035_ (.A(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .B(_06384_),
    .Y(_06438_));
 sky130_fd_sc_hd__o21ai_0 _25036_ (.A1(_10684_),
    .A2(_06437_),
    .B1(_06438_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _25037_ (.A(net3486),
    .B(_02990_),
    .Y(_06439_));
 sky130_fd_sc_hd__a21oi_1 _25038_ (.A1(net3683),
    .A2(_02990_),
    .B1(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _25039_ (.A(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .B(_06384_),
    .Y(_06441_));
 sky130_fd_sc_hd__o21ai_0 _25040_ (.A1(_10684_),
    .A2(_06440_),
    .B1(_06441_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _25041_ (.A(net3680),
    .B(net3631),
    .Y(_06442_));
 sky130_fd_sc_hd__a21oi_1 _25042_ (.A1(net168),
    .A2(net3631),
    .B1(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_114 ();
 sky130_fd_sc_hd__nand2_1 _25044_ (.A(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .B(_06384_),
    .Y(_06445_));
 sky130_fd_sc_hd__o21ai_0 _25045_ (.A1(_10684_),
    .A2(_06443_),
    .B1(_06445_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _25046_ (.A(_10294_),
    .B(net3631),
    .Y(_06446_));
 sky130_fd_sc_hd__a21oi_1 _25047_ (.A1(net169),
    .A2(net3631),
    .B1(_06446_),
    .Y(_06447_));
 sky130_fd_sc_hd__nand2_1 _25048_ (.A(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .B(_06384_),
    .Y(_06448_));
 sky130_fd_sc_hd__o21ai_0 _25049_ (.A1(_10684_),
    .A2(_06447_),
    .B1(_06448_),
    .Y(_01533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_113 ();
 sky130_fd_sc_hd__mux2i_1 _25051_ (.A0(net3474),
    .A1(_10360_),
    .S(_04421_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand2_1 _25052_ (.A(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .B(_06384_),
    .Y(_06451_));
 sky130_fd_sc_hd__o21ai_0 _25053_ (.A1(_10684_),
    .A2(_06450_),
    .B1(_06451_),
    .Y(_01534_));
 sky130_fd_sc_hd__mux2i_1 _25054_ (.A0(net3549),
    .A1(net3715),
    .S(_04421_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _25055_ (.A(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .B(_06384_),
    .Y(_06453_));
 sky130_fd_sc_hd__o21ai_0 _25056_ (.A1(_10684_),
    .A2(_06452_),
    .B1(_06453_),
    .Y(_01535_));
 sky130_fd_sc_hd__mux2i_1 _25057_ (.A0(net480),
    .A1(_10474_),
    .S(_04421_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand2_1 _25058_ (.A(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .B(_06384_),
    .Y(_06455_));
 sky130_fd_sc_hd__o21ai_0 _25059_ (.A1(_10684_),
    .A2(_06454_),
    .B1(_06455_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor3_1 _25060_ (.A(net471),
    .B(net3737),
    .C(net173),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_1 _25061_ (.A(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .B(_06384_),
    .Y(_06457_));
 sky130_fd_sc_hd__o31ai_1 _25062_ (.A1(_10390_),
    .A2(_10684_),
    .A3(_06456_),
    .B1(_06457_),
    .Y(_01537_));
 sky130_fd_sc_hd__or3_4 _25063_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(_07864_),
    .X(_06458_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_112 ();
 sky130_fd_sc_hd__nor2_4 _25065_ (.A(_13048_),
    .B(_06458_),
    .Y(_06460_));
 sky130_fd_sc_hd__a21oi_1 _25066_ (.A1(_13071_),
    .A2(_13189_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .Y(_06461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_111 ();
 sky130_fd_sc_hd__nand2_1 _25068_ (.A(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .B(_13181_),
    .Y(_06463_));
 sky130_fd_sc_hd__o21ai_2 _25069_ (.A1(net3575),
    .A2(_13181_),
    .B1(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__nor2_1 _25070_ (.A(_13048_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__a21oi_1 _25071_ (.A1(_13048_),
    .A2(_06461_),
    .B1(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__xnor2_1 _25072_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13071_),
    .Y(_06467_));
 sky130_fd_sc_hd__mux4_2 _25073_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06468_));
 sky130_fd_sc_hd__mux4_2 _25074_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_06469_));
 sky130_fd_sc_hd__mux4_2 _25075_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_06470_));
 sky130_fd_sc_hd__mux4_2 _25076_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_06471_));
 sky130_fd_sc_hd__mux4_2 _25077_ (.A0(_06468_),
    .A1(_06469_),
    .A2(_06470_),
    .A3(_06471_),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .X(_06472_));
 sky130_fd_sc_hd__a21oi_1 _25078_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B1(_10674_),
    .Y(_06473_));
 sky130_fd_sc_hd__mux2_1 _25079_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_06474_));
 sky130_fd_sc_hd__a21oi_1 _25080_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_06474_),
    .B1(_10672_),
    .Y(_06475_));
 sky130_fd_sc_hd__nor2_1 _25081_ (.A(_06473_),
    .B(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__o31ai_1 _25082_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B1(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__mux4_2 _25083_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06478_));
 sky130_fd_sc_hd__o22ai_1 _25084_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .A2(_13068_),
    .B1(_06476_),
    .B2(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__a21oi_1 _25085_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_06477_),
    .B1(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__mux4_2 _25086_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06481_));
 sky130_fd_sc_hd__mux4_2 _25087_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_06482_));
 sky130_fd_sc_hd__mux2i_1 _25088_ (.A0(_06481_),
    .A1(_06482_),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_06483_));
 sky130_fd_sc_hd__nor2_1 _25089_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__a21oi_2 _25090_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_06480_),
    .B1(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__nor2_1 _25091_ (.A(_06485_),
    .B(_06467_),
    .Y(_06486_));
 sky130_fd_sc_hd__a21oi_1 _25092_ (.A1(_06467_),
    .A2(_06472_),
    .B1(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nor3_4 _25093_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(_07864_),
    .Y(_06488_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__a21oi_1 _25095_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B1(_06488_),
    .Y(_06490_));
 sky130_fd_sc_hd__o221ai_1 _25096_ (.A1(_08169_),
    .A2(net3575),
    .B1(_06487_),
    .B2(_07862_),
    .C1(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__a21oi_2 _25097_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06466_),
    .B1(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__a211oi_1 _25099_ (.A1(net3711),
    .A2(_06460_),
    .B1(_06492_),
    .C1(_13047_),
    .Y(_06494_));
 sky130_fd_sc_hd__nor2_1 _25100_ (.A(_02225_),
    .B(_02977_),
    .Y(_06495_));
 sky130_fd_sc_hd__nor2_1 _25101_ (.A(_10690_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__o21ai_0 _25102_ (.A1(_13048_),
    .A2(_13098_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2_1 _25103_ (.A(_13078_),
    .B(_02990_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand3_1 _25104_ (.A(net3675),
    .B(_13048_),
    .C(net3631),
    .Y(_06499_));
 sky130_fd_sc_hd__a21oi_1 _25105_ (.A1(_06498_),
    .A2(_06499_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .Y(_06500_));
 sky130_fd_sc_hd__o22ai_1 _25106_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_06458_),
    .B1(_06497_),
    .B2(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_2 _25107_ (.A(net3937),
    .B(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand3_4 _25108_ (.A(net3755),
    .B(_10542_),
    .C(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__nor2_2 _25111_ (.A(_02225_),
    .B(_06503_),
    .Y(_06506_));
 sky130_fd_sc_hd__o32a_1 _25112_ (.A1(_06494_),
    .A2(_06496_),
    .A3(_06503_),
    .B1(_06506_),
    .B2(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .X(_01538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_103 ();
 sky130_fd_sc_hd__nand2_1 _25117_ (.A(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .B(_13181_),
    .Y(_06511_));
 sky130_fd_sc_hd__o21ai_0 _25118_ (.A1(_13118_),
    .A2(_13181_),
    .B1(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__or3_4 _25119_ (.A(net3940),
    .B(_08009_),
    .C(net3745),
    .X(_06513_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_102 ();
 sky130_fd_sc_hd__nor2_1 _25121_ (.A(_10676_),
    .B(_13181_),
    .Y(_06515_));
 sky130_fd_sc_hd__nor3_1 _25122_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .B(_06513_),
    .C(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nor2_1 _25123_ (.A(_07863_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__o21ai_0 _25124_ (.A1(_13048_),
    .A2(_06512_),
    .B1(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__a221oi_1 _25125_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3556),
    .B1(_06464_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_101 ();
 sky130_fd_sc_hd__nand2_4 _25127_ (.A(_06513_),
    .B(net3730),
    .Y(_06521_));
 sky130_fd_sc_hd__nor2_1 _25128_ (.A(net3714),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__a21oi_1 _25129_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__nor2_1 _25130_ (.A(_13047_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a31oi_1 _25131_ (.A1(_13047_),
    .A2(_02000_),
    .A3(_03104_),
    .B1(_06524_),
    .Y(_06525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_100 ();
 sky130_fd_sc_hd__o22a_1 _25133_ (.A1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A2(_06506_),
    .B1(_06525_),
    .B2(_06503_),
    .X(_01539_));
 sky130_fd_sc_hd__nor2_1 _25134_ (.A(_13192_),
    .B(_13240_),
    .Y(_06527_));
 sky130_fd_sc_hd__nor3_2 _25135_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .B(_06513_),
    .C(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_98 ();
 sky130_fd_sc_hd__nand2_1 _25138_ (.A(net171),
    .B(_13208_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _25139_ (.A(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B(_13181_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand2_1 _25140_ (.A(_06531_),
    .B(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__o21ai_0 _25141_ (.A1(_13048_),
    .A2(_06533_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06534_));
 sky130_fd_sc_hd__a221oi_1 _25142_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net171),
    .B1(_06512_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06535_));
 sky130_fd_sc_hd__o21ai_0 _25143_ (.A1(_06528_),
    .A2(_06534_),
    .B1(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__o21ai_2 _25144_ (.A1(net393),
    .A2(_06521_),
    .B1(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__nor3_1 _25145_ (.A(_10690_),
    .B(_02225_),
    .C(_03401_),
    .Y(_06538_));
 sky130_fd_sc_hd__a21oi_1 _25146_ (.A1(_10690_),
    .A2(_06537_),
    .B1(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__o22a_1 _25147_ (.A1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A2(_06506_),
    .B1(_06539_),
    .B2(_06503_),
    .X(_01540_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_97 ();
 sky130_fd_sc_hd__nor2_1 _25149_ (.A(_10690_),
    .B(_05069_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_1 _25150_ (.A(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B(_13181_),
    .Y(_06542_));
 sky130_fd_sc_hd__o21ai_2 _25151_ (.A1(net3534),
    .A2(_13181_),
    .B1(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__nor2_1 _25152_ (.A(_13195_),
    .B(_13240_),
    .Y(_06544_));
 sky130_fd_sc_hd__or3_4 _25153_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .B(_06513_),
    .C(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__o211ai_1 _25154_ (.A1(_13048_),
    .A2(_06543_),
    .B1(_06545_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__a221oi_1 _25156_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net174),
    .B1(_06533_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06548_));
 sky130_fd_sc_hd__o21ai_0 _25157_ (.A1(net3717),
    .A2(_06521_),
    .B1(net3734),
    .Y(_06549_));
 sky130_fd_sc_hd__a21oi_2 _25158_ (.A1(_06546_),
    .A2(_06548_),
    .B1(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__nor2_1 _25159_ (.A(_06541_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__nand2_1 _25161_ (.A(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B(_06503_),
    .Y(_06553_));
 sky130_fd_sc_hd__o21ai_0 _25162_ (.A1(_06503_),
    .A2(_06551_),
    .B1(_06553_),
    .Y(_01541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_93 ();
 sky130_fd_sc_hd__nand2_1 _25165_ (.A(net3536),
    .B(_13208_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand2_1 _25166_ (.A(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B(_13181_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_2 _25167_ (.A(_06556_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__a21oi_1 _25168_ (.A1(_13189_),
    .A2(_13219_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .Y(_06559_));
 sky130_fd_sc_hd__nand2_2 _25169_ (.A(_13048_),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__o211ai_1 _25170_ (.A1(_13048_),
    .A2(_06558_),
    .B1(_06560_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06561_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_91 ();
 sky130_fd_sc_hd__a221oi_1 _25173_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3536),
    .B1(_06543_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06564_));
 sky130_fd_sc_hd__a221oi_1 _25174_ (.A1(net3708),
    .A2(_06460_),
    .B1(_06561_),
    .B2(_06564_),
    .C1(_13047_),
    .Y(_06565_));
 sky130_fd_sc_hd__a21oi_1 _25175_ (.A1(_13047_),
    .A2(_03251_),
    .B1(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_1 _25176_ (.A(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B(_06503_),
    .Y(_06567_));
 sky130_fd_sc_hd__o21ai_0 _25177_ (.A1(_06503_),
    .A2(_06566_),
    .B1(_06567_),
    .Y(_01542_));
 sky130_fd_sc_hd__a221oi_1 _25178_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3537),
    .B1(_06558_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06568_));
 sky130_fd_sc_hd__or3_4 _25179_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13181_),
    .C(_13221_),
    .X(_06569_));
 sky130_fd_sc_hd__nor2_1 _25180_ (.A(_10674_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__mux2i_2 _25181_ (.A0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A1(net3537),
    .S(_13208_),
    .Y(_06571_));
 sky130_fd_sc_hd__a21oi_1 _25182_ (.A1(_06513_),
    .A2(_06571_),
    .B1(_07863_),
    .Y(_06572_));
 sky130_fd_sc_hd__o31ai_2 _25183_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .A2(_06513_),
    .A3(_06570_),
    .B1(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__a22oi_1 _25184_ (.A1(net376),
    .A2(_06460_),
    .B1(_06568_),
    .B2(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__nor2_1 _25185_ (.A(_13047_),
    .B(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__a31oi_1 _25186_ (.A1(_13047_),
    .A2(_02000_),
    .A3(_03764_),
    .B1(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__o22a_1 _25187_ (.A1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A2(_06506_),
    .B1(_06576_),
    .B2(_06503_),
    .X(_01543_));
 sky130_fd_sc_hd__nor2_1 _25188_ (.A(net3534),
    .B(_02990_),
    .Y(_06577_));
 sky130_fd_sc_hd__a21oi_1 _25189_ (.A1(net3719),
    .A2(_02990_),
    .B1(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__nand2_1 _25190_ (.A(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .B(_06384_),
    .Y(_06579_));
 sky130_fd_sc_hd__o21ai_0 _25191_ (.A1(_10684_),
    .A2(_06578_),
    .B1(_06579_),
    .Y(_01544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_89 ();
 sky130_fd_sc_hd__nor2_1 _25194_ (.A(net3529),
    .B(_13181_),
    .Y(_06582_));
 sky130_fd_sc_hd__a21oi_2 _25195_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_13181_),
    .B1(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__a211oi_2 _25196_ (.A1(_13057_),
    .A2(_01646_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .C1(_06513_),
    .Y(_06584_));
 sky130_fd_sc_hd__a21oi_1 _25197_ (.A1(_06513_),
    .A2(_06583_),
    .B1(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__o221ai_1 _25198_ (.A1(_08169_),
    .A2(net3529),
    .B1(_06571_),
    .B2(_07862_),
    .C1(_06458_),
    .Y(_06586_));
 sky130_fd_sc_hd__a21oi_2 _25199_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06585_),
    .B1(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__a21oi_1 _25200_ (.A1(net3724),
    .A2(_06460_),
    .B1(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_88 ();
 sky130_fd_sc_hd__nor2_1 _25202_ (.A(_10690_),
    .B(_04936_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_1 _25203_ (.A1(_10690_),
    .A2(_06588_),
    .B1(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _25204_ (.A(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .B(_06503_),
    .Y(_06592_));
 sky130_fd_sc_hd__o21ai_0 _25205_ (.A1(_06503_),
    .A2(_06591_),
    .B1(_06592_),
    .Y(_01545_));
 sky130_fd_sc_hd__nor2_1 _25206_ (.A(_13195_),
    .B(_06569_),
    .Y(_06593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_87 ();
 sky130_fd_sc_hd__mux2i_1 _25208_ (.A0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A1(net3530),
    .S(_13208_),
    .Y(_06595_));
 sky130_fd_sc_hd__nand2_1 _25209_ (.A(_06513_),
    .B(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_86 ();
 sky130_fd_sc_hd__o311ai_0 _25211_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .A2(_06513_),
    .A3(_06593_),
    .B1(_06596_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06598_));
 sky130_fd_sc_hd__a21oi_1 _25212_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3530),
    .B1(_06488_),
    .Y(_06599_));
 sky130_fd_sc_hd__o211ai_1 _25213_ (.A1(_07862_),
    .A2(_06583_),
    .B1(_06598_),
    .C1(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__a21oi_1 _25214_ (.A1(net403),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06601_));
 sky130_fd_sc_hd__a22oi_1 _25215_ (.A1(_13047_),
    .A2(_04952_),
    .B1(_06600_),
    .B2(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__nand2_1 _25216_ (.A(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B(_06503_),
    .Y(_06603_));
 sky130_fd_sc_hd__o21ai_0 _25217_ (.A1(_06503_),
    .A2(_06602_),
    .B1(_06603_),
    .Y(_01546_));
 sky130_fd_sc_hd__mux2i_1 _25218_ (.A0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .A1(net3519),
    .S(_13208_),
    .Y(_06604_));
 sky130_fd_sc_hd__a211oi_2 _25219_ (.A1(_13067_),
    .A2(_13199_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .C1(_06513_),
    .Y(_06605_));
 sky130_fd_sc_hd__a21oi_1 _25220_ (.A1(_06513_),
    .A2(_06604_),
    .B1(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__a21oi_1 _25221_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3519),
    .B1(_06488_),
    .Y(_06607_));
 sky130_fd_sc_hd__o21ai_0 _25222_ (.A1(_07862_),
    .A2(_06595_),
    .B1(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__a21oi_1 _25223_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06606_),
    .B1(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__o21ai_0 _25224_ (.A1(net3704),
    .A2(_06521_),
    .B1(net3734),
    .Y(_06610_));
 sky130_fd_sc_hd__o22a_1 _25225_ (.A1(net3734),
    .A2(_02003_),
    .B1(_06609_),
    .B2(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__nand2_1 _25226_ (.A(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .B(_06503_),
    .Y(_06612_));
 sky130_fd_sc_hd__o21ai_0 _25227_ (.A1(_06503_),
    .A2(_06611_),
    .B1(_06612_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand2_1 _25228_ (.A(net3520),
    .B(_13208_),
    .Y(_06613_));
 sky130_fd_sc_hd__nand2_1 _25229_ (.A(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B(_13181_),
    .Y(_06614_));
 sky130_fd_sc_hd__nand2_1 _25230_ (.A(_06613_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__o21ai_0 _25231_ (.A1(_13048_),
    .A2(_06615_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06616_));
 sky130_fd_sc_hd__a311oi_1 _25232_ (.A1(_10672_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13191_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .Y(_06617_));
 sky130_fd_sc_hd__a21oi_1 _25233_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3520),
    .B1(_06488_),
    .Y(_06618_));
 sky130_fd_sc_hd__o221ai_1 _25234_ (.A1(_07862_),
    .A2(_06604_),
    .B1(_06616_),
    .B2(_06617_),
    .C1(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__a21oi_1 _25235_ (.A1(net3705),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06620_));
 sky130_fd_sc_hd__nor2_1 _25236_ (.A(_10690_),
    .B(_02291_),
    .Y(_06621_));
 sky130_fd_sc_hd__a21oi_1 _25237_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_85 ();
 sky130_fd_sc_hd__nand2_1 _25239_ (.A(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B(_06503_),
    .Y(_06624_));
 sky130_fd_sc_hd__o21ai_0 _25240_ (.A1(_06503_),
    .A2(_06622_),
    .B1(_06624_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _25241_ (.A(net151),
    .B(_13208_),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_1 _25242_ (.A(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B(_13181_),
    .Y(_06626_));
 sky130_fd_sc_hd__nand2_1 _25243_ (.A(_06625_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21ai_0 _25244_ (.A1(_13048_),
    .A2(_06627_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06628_));
 sky130_fd_sc_hd__a211oi_2 _25245_ (.A1(_13057_),
    .A2(_13191_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .C1(_06513_),
    .Y(_06629_));
 sky130_fd_sc_hd__a221oi_1 _25246_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net151),
    .B1(_06615_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06630_));
 sky130_fd_sc_hd__o21ai_2 _25247_ (.A1(_06628_),
    .A2(_06629_),
    .B1(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__a21oi_1 _25248_ (.A1(net400),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06632_));
 sky130_fd_sc_hd__nor2_1 _25249_ (.A(_10690_),
    .B(_02385_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21oi_1 _25250_ (.A1(_06631_),
    .A2(_06632_),
    .B1(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__nand2_1 _25251_ (.A(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B(_06503_),
    .Y(_06635_));
 sky130_fd_sc_hd__o21ai_0 _25252_ (.A1(_06503_),
    .A2(_06634_),
    .B1(_06635_),
    .Y(_01549_));
 sky130_fd_sc_hd__nand2_1 _25253_ (.A(net152),
    .B(_13208_),
    .Y(_06636_));
 sky130_fd_sc_hd__nand2_1 _25254_ (.A(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B(_13181_),
    .Y(_06637_));
 sky130_fd_sc_hd__nand2_1 _25255_ (.A(_06636_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__o21ai_0 _25256_ (.A1(_13048_),
    .A2(_06638_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06639_));
 sky130_fd_sc_hd__a311oi_2 _25257_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13191_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .Y(_06640_));
 sky130_fd_sc_hd__a221oi_1 _25258_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net152),
    .B1(_06627_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06641_));
 sky130_fd_sc_hd__o21ai_0 _25259_ (.A1(_06639_),
    .A2(_06640_),
    .B1(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21oi_1 _25260_ (.A1(net3703),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06643_));
 sky130_fd_sc_hd__nor2_1 _25261_ (.A(net3734),
    .B(_02531_),
    .Y(_06644_));
 sky130_fd_sc_hd__a21oi_1 _25262_ (.A1(_06642_),
    .A2(_06643_),
    .B1(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand2_1 _25263_ (.A(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B(_06503_),
    .Y(_06646_));
 sky130_fd_sc_hd__o21ai_0 _25264_ (.A1(_06503_),
    .A2(_06645_),
    .B1(_06646_),
    .Y(_01550_));
 sky130_fd_sc_hd__inv_1 _25265_ (.A(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .Y(_06647_));
 sky130_fd_sc_hd__nor2_1 _25266_ (.A(net3734),
    .B(_02606_),
    .Y(_06648_));
 sky130_fd_sc_hd__nor2_1 _25267_ (.A(_13218_),
    .B(_13190_),
    .Y(_06649_));
 sky130_fd_sc_hd__mux2i_1 _25268_ (.A0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A1(net3514),
    .S(_13208_),
    .Y(_06650_));
 sky130_fd_sc_hd__nand2_1 _25269_ (.A(_06513_),
    .B(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__o311ai_1 _25270_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .A2(_06513_),
    .A3(_06649_),
    .B1(_06651_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06652_));
 sky130_fd_sc_hd__a221oi_1 _25271_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3514),
    .B1(_06638_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06653_));
 sky130_fd_sc_hd__a221oi_1 _25272_ (.A1(net401),
    .A2(_06460_),
    .B1(_06652_),
    .B2(_06653_),
    .C1(_13047_),
    .Y(_06654_));
 sky130_fd_sc_hd__nor3_1 _25273_ (.A(_06503_),
    .B(_06648_),
    .C(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__a21oi_1 _25274_ (.A1(_06647_),
    .A2(_06503_),
    .B1(_06655_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _25275_ (.A(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B(_13181_),
    .Y(_06656_));
 sky130_fd_sc_hd__o21ai_2 _25276_ (.A1(net3498),
    .A2(_13181_),
    .B1(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__o21ai_0 _25277_ (.A1(_13048_),
    .A2(_06657_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06658_));
 sky130_fd_sc_hd__a311oi_1 _25278_ (.A1(_10672_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13201_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .Y(_06659_));
 sky130_fd_sc_hd__a21oi_1 _25279_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net154),
    .B1(_06488_),
    .Y(_06660_));
 sky130_fd_sc_hd__o221ai_1 _25280_ (.A1(_07862_),
    .A2(_06650_),
    .B1(_06658_),
    .B2(_06659_),
    .C1(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__a21oi_1 _25281_ (.A1(net3699),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06662_));
 sky130_fd_sc_hd__nor2_1 _25282_ (.A(net3734),
    .B(_02699_),
    .Y(_06663_));
 sky130_fd_sc_hd__a21oi_1 _25283_ (.A1(_06661_),
    .A2(_06662_),
    .B1(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_1 _25284_ (.A(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B(_06503_),
    .Y(_06665_));
 sky130_fd_sc_hd__o21ai_0 _25285_ (.A1(_06503_),
    .A2(_06664_),
    .B1(_06665_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _25286_ (.A(net3734),
    .B(_06503_),
    .Y(_06666_));
 sky130_fd_sc_hd__a21oi_2 _25287_ (.A1(_13057_),
    .A2(_13201_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2_1 _25288_ (.A(net3513),
    .B(_13208_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_1 _25289_ (.A(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B(_13181_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand2_1 _25290_ (.A(_06668_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__nor2_1 _25291_ (.A(_13048_),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__a21oi_1 _25292_ (.A1(_13048_),
    .A2(_06667_),
    .B1(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__a221o_1 _25293_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3513),
    .B1(_06657_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .X(_06673_));
 sky130_fd_sc_hd__a21oi_1 _25294_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06672_),
    .B1(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__a2111oi_0 _25295_ (.A1(net3695),
    .A2(_06460_),
    .B1(_06503_),
    .C1(_06674_),
    .D1(_13047_),
    .Y(_06675_));
 sky130_fd_sc_hd__a221o_1 _25296_ (.A1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A2(_06503_),
    .B1(_06666_),
    .B2(_02816_),
    .C1(_06675_),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _25297_ (.A(net3507),
    .B(_13208_),
    .Y(_06676_));
 sky130_fd_sc_hd__nand2_1 _25298_ (.A(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B(_13181_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_1 _25299_ (.A(_06676_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21ai_0 _25300_ (.A1(_13048_),
    .A2(_06678_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06679_));
 sky130_fd_sc_hd__a311oi_2 _25301_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13201_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .Y(_06680_));
 sky130_fd_sc_hd__a221oi_1 _25302_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3507),
    .B1(_06670_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06681_));
 sky130_fd_sc_hd__o21ai_0 _25303_ (.A1(_06679_),
    .A2(_06680_),
    .B1(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__a21oi_1 _25304_ (.A1(net3697),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06683_));
 sky130_fd_sc_hd__nor2_1 _25305_ (.A(net3734),
    .B(_02944_),
    .Y(_06684_));
 sky130_fd_sc_hd__a21oi_1 _25306_ (.A1(_06682_),
    .A2(_06683_),
    .B1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand2_1 _25307_ (.A(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B(_06503_),
    .Y(_06686_));
 sky130_fd_sc_hd__o21ai_0 _25308_ (.A1(_06503_),
    .A2(_06685_),
    .B1(_06686_),
    .Y(_01554_));
 sky130_fd_sc_hd__mux2i_1 _25309_ (.A0(net3707),
    .A1(net3536),
    .S(net3631),
    .Y(_06687_));
 sky130_fd_sc_hd__nand2_1 _25310_ (.A(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .B(_06384_),
    .Y(_06688_));
 sky130_fd_sc_hd__o21ai_0 _25311_ (.A1(_10684_),
    .A2(_06687_),
    .B1(_06688_),
    .Y(_01555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_84 ();
 sky130_fd_sc_hd__mux2i_1 _25313_ (.A0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .A1(net3506),
    .S(_13208_),
    .Y(_06690_));
 sky130_fd_sc_hd__a211oi_1 _25314_ (.A1(_13071_),
    .A2(_13229_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .C1(_06513_),
    .Y(_06691_));
 sky130_fd_sc_hd__a21oi_1 _25315_ (.A1(_06513_),
    .A2(_06690_),
    .B1(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a221o_1 _25316_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3506),
    .B1(_06678_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .X(_06693_));
 sky130_fd_sc_hd__a21oi_1 _25317_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06692_),
    .B1(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__a21oi_1 _25318_ (.A1(net3693),
    .A2(_06460_),
    .B1(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__nor2_1 _25319_ (.A(net3734),
    .B(_03081_),
    .Y(_06696_));
 sky130_fd_sc_hd__a21oi_1 _25320_ (.A1(net3734),
    .A2(_06695_),
    .B1(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_1 _25321_ (.A(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B(_06503_),
    .Y(_06698_));
 sky130_fd_sc_hd__o21ai_0 _25322_ (.A1(_06503_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand2_1 _25323_ (.A(net420),
    .B(_13208_),
    .Y(_06699_));
 sky130_fd_sc_hd__nand2_1 _25324_ (.A(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B(_13181_),
    .Y(_06700_));
 sky130_fd_sc_hd__nand2_1 _25325_ (.A(_06699_),
    .B(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nor2_1 _25326_ (.A(_13048_),
    .B(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__a211oi_1 _25327_ (.A1(_10675_),
    .A2(_13229_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .Y(_06703_));
 sky130_fd_sc_hd__nor3_1 _25328_ (.A(_07863_),
    .B(_06702_),
    .C(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__nor2_1 _25329_ (.A(_07862_),
    .B(_06690_),
    .Y(_06705_));
 sky130_fd_sc_hd__a2111oi_1 _25330_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net420),
    .B1(_06488_),
    .C1(_06704_),
    .D1(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__o21ai_0 _25331_ (.A1(net332),
    .A2(_06521_),
    .B1(net3734),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_1 _25332_ (.A(_13047_),
    .B(_03218_),
    .Y(_06708_));
 sky130_fd_sc_hd__o21ai_0 _25333_ (.A1(_06706_),
    .A2(_06707_),
    .B1(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__mux2_1 _25334_ (.A0(_06709_),
    .A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .S(_06503_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _25335_ (.A(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B(_13181_),
    .Y(_06710_));
 sky130_fd_sc_hd__o21ai_0 _25336_ (.A1(net3497),
    .A2(_13181_),
    .B1(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__o21ai_0 _25337_ (.A1(_13048_),
    .A2(_06711_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06712_));
 sky130_fd_sc_hd__a211oi_2 _25338_ (.A1(_13057_),
    .A2(_13213_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .C1(_06513_),
    .Y(_06713_));
 sky130_fd_sc_hd__a221oi_1 _25339_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net159),
    .B1(_06701_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06714_));
 sky130_fd_sc_hd__o21ai_0 _25340_ (.A1(_06712_),
    .A2(_06713_),
    .B1(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__a21oi_1 _25341_ (.A1(_09652_),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06716_));
 sky130_fd_sc_hd__a22oi_1 _25342_ (.A1(_13047_),
    .A2(_03403_),
    .B1(_06715_),
    .B2(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_1 _25343_ (.A(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B(_06503_),
    .Y(_06718_));
 sky130_fd_sc_hd__o21ai_0 _25344_ (.A1(_06503_),
    .A2(_06717_),
    .B1(_06718_),
    .Y(_01558_));
 sky130_fd_sc_hd__a31oi_2 _25345_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13213_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_1 _25346_ (.A(net160),
    .B(_13208_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand2_1 _25347_ (.A(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B(_13181_),
    .Y(_06721_));
 sky130_fd_sc_hd__nand2_1 _25348_ (.A(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__nor2_1 _25349_ (.A(_13048_),
    .B(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21oi_1 _25350_ (.A1(_13048_),
    .A2(_06719_),
    .B1(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__a221o_1 _25351_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net160),
    .B1(_06711_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .X(_06725_));
 sky130_fd_sc_hd__a21oi_1 _25352_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06724_),
    .B1(_06725_),
    .Y(_06726_));
 sky130_fd_sc_hd__o21ai_0 _25353_ (.A1(net422),
    .A2(_06521_),
    .B1(net3734),
    .Y(_06727_));
 sky130_fd_sc_hd__nor2_1 _25354_ (.A(_06726_),
    .B(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__a21oi_1 _25355_ (.A1(_13047_),
    .A2(_03519_),
    .B1(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_1 _25356_ (.A(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B(_06503_),
    .Y(_06730_));
 sky130_fd_sc_hd__o21ai_0 _25357_ (.A1(_06503_),
    .A2(_06729_),
    .B1(_06730_),
    .Y(_01559_));
 sky130_fd_sc_hd__mux2i_1 _25358_ (.A0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A1(net452),
    .S(_13208_),
    .Y(_06731_));
 sky130_fd_sc_hd__a211oi_2 _25359_ (.A1(_13229_),
    .A2(_13219_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .C1(_06513_),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_1 _25360_ (.A1(_06513_),
    .A2(_06731_),
    .B1(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_1 _25361_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__a221oi_1 _25362_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net452),
    .B1(_06722_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(net3730),
    .Y(_06735_));
 sky130_fd_sc_hd__a221oi_2 _25363_ (.A1(net3689),
    .A2(_06460_),
    .B1(_06734_),
    .B2(_06735_),
    .C1(_13047_),
    .Y(_06736_));
 sky130_fd_sc_hd__a21oi_1 _25364_ (.A1(_13047_),
    .A2(_03642_),
    .B1(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_1 _25365_ (.A(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .B(_06503_),
    .Y(_06738_));
 sky130_fd_sc_hd__o21ai_0 _25366_ (.A1(_06503_),
    .A2(_06737_),
    .B1(_06738_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _25367_ (.A(net3496),
    .B(_13181_),
    .Y(_06739_));
 sky130_fd_sc_hd__a21oi_1 _25368_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_13181_),
    .B1(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__nand2_1 _25369_ (.A(_06513_),
    .B(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__a311o_1 _25370_ (.A1(_10672_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13222_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .X(_06742_));
 sky130_fd_sc_hd__nor2_1 _25371_ (.A(_07862_),
    .B(_06731_),
    .Y(_06743_));
 sky130_fd_sc_hd__o21ai_0 _25372_ (.A1(_08169_),
    .A2(net3496),
    .B1(_06458_),
    .Y(_06744_));
 sky130_fd_sc_hd__a311o_1 _25373_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06741_),
    .A3(_06742_),
    .B1(_06743_),
    .C1(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__a21oi_1 _25374_ (.A1(net3690),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06746_));
 sky130_fd_sc_hd__a21oi_1 _25375_ (.A1(_02000_),
    .A2(_03760_),
    .B1(_03765_),
    .Y(_06747_));
 sky130_fd_sc_hd__nor2_1 _25376_ (.A(_10690_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__a21oi_1 _25377_ (.A1(_06745_),
    .A2(_06746_),
    .B1(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _25378_ (.A(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B(_06503_),
    .Y(_06750_));
 sky130_fd_sc_hd__o21ai_0 _25379_ (.A1(_06503_),
    .A2(_06749_),
    .B1(_06750_),
    .Y(_01561_));
 sky130_fd_sc_hd__mux2i_1 _25380_ (.A0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A1(net3503),
    .S(_13208_),
    .Y(_06751_));
 sky130_fd_sc_hd__nor2_1 _25381_ (.A(_13048_),
    .B(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__a21oi_1 _25382_ (.A1(_13057_),
    .A2(_13222_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .Y(_06753_));
 sky130_fd_sc_hd__nor2_1 _25383_ (.A(_06513_),
    .B(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__o21ai_0 _25384_ (.A1(_06752_),
    .A2(_06754_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06755_));
 sky130_fd_sc_hd__a21oi_1 _25385_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3503),
    .B1(net3730),
    .Y(_06756_));
 sky130_fd_sc_hd__o21a_1 _25386_ (.A1(_07862_),
    .A2(_06740_),
    .B1(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__a221oi_2 _25387_ (.A1(net3687),
    .A2(_06460_),
    .B1(_06755_),
    .B2(_06757_),
    .C1(_13047_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21oi_1 _25388_ (.A1(_13047_),
    .A2(_03887_),
    .B1(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _25389_ (.A(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .B(_06503_),
    .Y(_06760_));
 sky130_fd_sc_hd__o21ai_0 _25390_ (.A1(_06503_),
    .A2(_06759_),
    .B1(_06760_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _25391_ (.A(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B(_13181_),
    .Y(_06761_));
 sky130_fd_sc_hd__o21ai_0 _25392_ (.A1(net3504),
    .A2(_13181_),
    .B1(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__a311o_1 _25393_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13222_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .X(_06763_));
 sky130_fd_sc_hd__o211ai_1 _25394_ (.A1(_13048_),
    .A2(_06762_),
    .B1(_06763_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06764_));
 sky130_fd_sc_hd__o221a_1 _25395_ (.A1(_08169_),
    .A2(net3504),
    .B1(_06751_),
    .B2(_07862_),
    .C1(_06458_),
    .X(_06765_));
 sky130_fd_sc_hd__a221oi_1 _25396_ (.A1(_09903_),
    .A2(_06460_),
    .B1(_06764_),
    .B2(_06765_),
    .C1(_13047_),
    .Y(_06766_));
 sky130_fd_sc_hd__o21ai_4 _25397_ (.A1(_03904_),
    .A2(net3432),
    .B1(_13047_),
    .Y(_06767_));
 sky130_fd_sc_hd__nor2b_1 _25398_ (.A(_06766_),
    .B_N(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand2_1 _25399_ (.A(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B(_06503_),
    .Y(_06769_));
 sky130_fd_sc_hd__o21ai_0 _25400_ (.A1(_06503_),
    .A2(_06768_),
    .B1(_06769_),
    .Y(_01563_));
 sky130_fd_sc_hd__mux2i_1 _25401_ (.A0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A1(net272),
    .S(_13208_),
    .Y(_06770_));
 sky130_fd_sc_hd__nor2_1 _25402_ (.A(_13048_),
    .B(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21oi_1 _25403_ (.A1(_13067_),
    .A2(_13226_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .Y(_06772_));
 sky130_fd_sc_hd__nor2_1 _25404_ (.A(_06513_),
    .B(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__o21ai_0 _25405_ (.A1(_06771_),
    .A2(_06773_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06774_));
 sky130_fd_sc_hd__a221oi_1 _25406_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net272),
    .B1(_06762_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06775_));
 sky130_fd_sc_hd__a221oi_1 _25407_ (.A1(_09983_),
    .A2(_06460_),
    .B1(_06774_),
    .B2(_06775_),
    .C1(_13047_),
    .Y(_06776_));
 sky130_fd_sc_hd__a21oi_1 _25408_ (.A1(_13047_),
    .A2(net3431),
    .B1(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_1 _25409_ (.A(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .B(_06503_),
    .Y(_06778_));
 sky130_fd_sc_hd__o21ai_0 _25410_ (.A1(_06503_),
    .A2(_06777_),
    .B1(_06778_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _25411_ (.A(_07862_),
    .B(_06770_),
    .Y(_06779_));
 sky130_fd_sc_hd__a211oi_1 _25412_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net3495),
    .B1(_06488_),
    .C1(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__mux2i_1 _25413_ (.A0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A1(net3495),
    .S(_13208_),
    .Y(_06781_));
 sky130_fd_sc_hd__nand2_1 _25414_ (.A(_06513_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__a311o_1 _25415_ (.A1(_10672_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A3(_13231_),
    .B1(_06513_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .X(_06783_));
 sky130_fd_sc_hd__nand3_1 _25416_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_06782_),
    .C(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__a221oi_2 _25417_ (.A1(_10088_),
    .A2(_06460_),
    .B1(_06780_),
    .B2(_06784_),
    .C1(_13047_),
    .Y(_06785_));
 sky130_fd_sc_hd__a21oi_1 _25418_ (.A1(_13047_),
    .A2(net3424),
    .B1(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__nand2_1 _25419_ (.A(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .B(_06503_),
    .Y(_06787_));
 sky130_fd_sc_hd__o21ai_0 _25420_ (.A1(_06503_),
    .A2(_06786_),
    .B1(_06787_),
    .Y(_01565_));
 sky130_fd_sc_hd__mux2i_1 _25421_ (.A0(net3537),
    .A1(_08240_),
    .S(_04421_),
    .Y(_06788_));
 sky130_fd_sc_hd__nand2_1 _25422_ (.A(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .B(_06384_),
    .Y(_06789_));
 sky130_fd_sc_hd__o21ai_0 _25423_ (.A1(_10684_),
    .A2(_06788_),
    .B1(_06789_),
    .Y(_01566_));
 sky130_fd_sc_hd__a21oi_1 _25424_ (.A1(_13057_),
    .A2(_13231_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .Y(_06790_));
 sky130_fd_sc_hd__nand2_1 _25425_ (.A(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .B(_13181_),
    .Y(_06791_));
 sky130_fd_sc_hd__o21ai_0 _25426_ (.A1(net3486),
    .A2(_13181_),
    .B1(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__nor2_1 _25427_ (.A(_13048_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21oi_2 _25428_ (.A1(_13048_),
    .A2(_06790_),
    .B1(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__o221ai_1 _25429_ (.A1(_08169_),
    .A2(net3486),
    .B1(_06781_),
    .B2(_07862_),
    .C1(_06458_),
    .Y(_06795_));
 sky130_fd_sc_hd__a21oi_4 _25430_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06794_),
    .B1(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__a2111oi_0 _25431_ (.A1(net3682),
    .A2(_06460_),
    .B1(_06503_),
    .C1(_06796_),
    .D1(_13047_),
    .Y(_06797_));
 sky130_fd_sc_hd__nor4_2 _25432_ (.A(_10690_),
    .B(_04250_),
    .C(_04349_),
    .D(_06503_),
    .Y(_06798_));
 sky130_fd_sc_hd__a211o_1 _25433_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_06503_),
    .B1(_06797_),
    .C1(_06798_),
    .X(_01567_));
 sky130_fd_sc_hd__a221oi_1 _25434_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net168),
    .B1(_06792_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06799_));
 sky130_fd_sc_hd__nor3_1 _25435_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13195_),
    .C(_13230_),
    .Y(_06800_));
 sky130_fd_sc_hd__nor2_1 _25436_ (.A(net3487),
    .B(_13181_),
    .Y(_06801_));
 sky130_fd_sc_hd__a21oi_2 _25437_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(_13181_),
    .B1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand2_1 _25438_ (.A(_06513_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__o311ai_2 _25439_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .A2(_06513_),
    .A3(_06800_),
    .B1(_06803_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06804_));
 sky130_fd_sc_hd__a221oi_4 _25440_ (.A1(net3681),
    .A2(_06460_),
    .B1(_06799_),
    .B2(_06804_),
    .C1(_13047_),
    .Y(_06805_));
 sky130_fd_sc_hd__a21oi_1 _25441_ (.A1(_04374_),
    .A2(_04447_),
    .B1(_10690_),
    .Y(_06806_));
 sky130_fd_sc_hd__nor3_1 _25442_ (.A(_06503_),
    .B(_06805_),
    .C(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__a21oi_1 _25443_ (.A1(_10204_),
    .A2(_06503_),
    .B1(_06807_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _25444_ (.A(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B(_13181_),
    .Y(_06808_));
 sky130_fd_sc_hd__o21ai_0 _25445_ (.A1(net3485),
    .A2(_13181_),
    .B1(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__a21oi_1 _25446_ (.A1(_13063_),
    .A2(_13226_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .Y(_06810_));
 sky130_fd_sc_hd__nor2_1 _25447_ (.A(_06513_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__a21oi_1 _25448_ (.A1(_06513_),
    .A2(_06809_),
    .B1(_06811_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21oi_1 _25449_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net169),
    .B1(_06488_),
    .Y(_06813_));
 sky130_fd_sc_hd__o221ai_2 _25450_ (.A1(_07862_),
    .A2(_06802_),
    .B1(_06812_),
    .B2(_07863_),
    .C1(_06813_),
    .Y(_06814_));
 sky130_fd_sc_hd__a21oi_1 _25451_ (.A1(net3679),
    .A2(_06460_),
    .B1(_13047_),
    .Y(_06815_));
 sky130_fd_sc_hd__nor2_1 _25452_ (.A(_10690_),
    .B(_04565_),
    .Y(_06816_));
 sky130_fd_sc_hd__a21oi_1 _25453_ (.A1(_06814_),
    .A2(_06815_),
    .B1(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_1 _25454_ (.A(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B(_06503_),
    .Y(_06818_));
 sky130_fd_sc_hd__o21ai_0 _25455_ (.A1(_06503_),
    .A2(_06817_),
    .B1(_06818_),
    .Y(_01569_));
 sky130_fd_sc_hd__a21oi_1 _25456_ (.A1(_02000_),
    .A2(net3423),
    .B1(_04677_),
    .Y(_06819_));
 sky130_fd_sc_hd__nand2_1 _25457_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13226_),
    .Y(_06820_));
 sky130_fd_sc_hd__nor2_1 _25458_ (.A(_10674_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__mux2i_1 _25459_ (.A0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A1(net292),
    .S(_13208_),
    .Y(_06822_));
 sky130_fd_sc_hd__nand2_1 _25460_ (.A(_06513_),
    .B(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__o311ai_1 _25461_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .A2(_06513_),
    .A3(_06821_),
    .B1(_06823_),
    .C1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06824_));
 sky130_fd_sc_hd__a221oi_1 _25462_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net292),
    .B1(_06809_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06825_));
 sky130_fd_sc_hd__a221oi_2 _25463_ (.A1(net3676),
    .A2(_06460_),
    .B1(_06824_),
    .B2(_06825_),
    .C1(_13047_),
    .Y(_06826_));
 sky130_fd_sc_hd__a21oi_1 _25464_ (.A1(_13047_),
    .A2(_06819_),
    .B1(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__nand2_1 _25465_ (.A(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .B(_06503_),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_0 _25466_ (.A1(_06503_),
    .A2(_06827_),
    .B1(_06828_),
    .Y(_01570_));
 sky130_fd_sc_hd__a21oi_1 _25467_ (.A1(_13057_),
    .A2(_13237_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_1 _25468_ (.A(net481),
    .B(_13208_),
    .Y(_06830_));
 sky130_fd_sc_hd__nand2_1 _25469_ (.A(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B(_13181_),
    .Y(_06831_));
 sky130_fd_sc_hd__nand2_1 _25470_ (.A(_06830_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nor2_1 _25471_ (.A(_13048_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__a21oi_1 _25472_ (.A1(_13048_),
    .A2(_06829_),
    .B1(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__a21oi_1 _25473_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net481),
    .B1(_06488_),
    .Y(_06835_));
 sky130_fd_sc_hd__o21ai_0 _25474_ (.A1(_07862_),
    .A2(_06822_),
    .B1(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(net3674),
    .B(_06460_),
    .Y(_06837_));
 sky130_fd_sc_hd__a22oi_1 _25476_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06834_),
    .B1(_06836_),
    .B2(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_1 _25477_ (.A(_13047_),
    .B(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__a21oi_1 _25478_ (.A1(_13047_),
    .A2(net3429),
    .B1(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand2_1 _25479_ (.A(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B(_06503_),
    .Y(_06841_));
 sky130_fd_sc_hd__o21ai_0 _25480_ (.A1(_06503_),
    .A2(_06840_),
    .B1(_06841_),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _25481_ (.A(_02225_),
    .B(_02942_),
    .Y(_06842_));
 sky130_fd_sc_hd__a21oi_2 _25482_ (.A1(net3422),
    .A2(_06842_),
    .B1(_10690_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_1 _25483_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .B(_13048_),
    .Y(_06844_));
 sky130_fd_sc_hd__nand3_1 _25484_ (.A(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B(net173),
    .C(_06513_),
    .Y(_06845_));
 sky130_fd_sc_hd__o311ai_0 _25485_ (.A1(net3940),
    .A2(_13195_),
    .A3(_06820_),
    .B1(_06844_),
    .C1(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a221oi_1 _25486_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net173),
    .B1(_06832_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06488_),
    .Y(_06847_));
 sky130_fd_sc_hd__a21oi_1 _25487_ (.A1(net3675),
    .A2(_06460_),
    .B1(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__a211oi_1 _25488_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06846_),
    .B1(_06848_),
    .C1(_13047_),
    .Y(_06849_));
 sky130_fd_sc_hd__nand2_1 _25489_ (.A(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B(_06503_),
    .Y(_06850_));
 sky130_fd_sc_hd__o31ai_1 _25490_ (.A1(_06503_),
    .A2(_06843_),
    .A3(_06849_),
    .B1(_06850_),
    .Y(_01572_));
 sky130_fd_sc_hd__o21ai_2 _25491_ (.A1(net3940),
    .A2(_06458_),
    .B1(net3734),
    .Y(_06851_));
 sky130_fd_sc_hd__a31oi_1 _25492_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A3(net173),
    .B1(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2b_1 _25493_ (.A_N(_04882_),
    .B(_04883_),
    .Y(_06853_));
 sky130_fd_sc_hd__inv_1 _25494_ (.A(_04807_),
    .Y(_06854_));
 sky130_fd_sc_hd__nor2_1 _25495_ (.A(net3450),
    .B(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nand2_1 _25496_ (.A(net3450),
    .B(_06854_),
    .Y(_06856_));
 sky130_fd_sc_hd__o21ai_0 _25497_ (.A1(_04732_),
    .A2(_06855_),
    .B1(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2b_2 _25498_ (.A(_04883_),
    .B_N(_04882_),
    .Y(_06858_));
 sky130_fd_sc_hd__a21oi_1 _25499_ (.A1(_06853_),
    .A2(_06857_),
    .B1(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__maj3_1 _25500_ (.A(_04819_),
    .B(_04877_),
    .C(_04881_),
    .X(_06860_));
 sky130_fd_sc_hd__nor2_1 _25501_ (.A(_04835_),
    .B(_04845_),
    .Y(_06861_));
 sky130_fd_sc_hd__nor2_1 _25502_ (.A(_04747_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21o_4 _25503_ (.A1(_04835_),
    .A2(_04845_),
    .B1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__nor2_1 _25504_ (.A(_04847_),
    .B(_04875_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand2_1 _25505_ (.A(_04847_),
    .B(_04875_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_2 _25506_ (.A1(_04834_),
    .A2(_06864_),
    .B1(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__a21o_4 _25507_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net3668),
    .B1(net3732),
    .X(_06867_));
 sky130_fd_sc_hd__nor2_1 _25508_ (.A(_04820_),
    .B(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__nor3_1 _25509_ (.A(_03460_),
    .B(_03803_),
    .C(_06867_),
    .Y(_06869_));
 sky130_fd_sc_hd__a311oi_1 _25510_ (.A1(_03460_),
    .A2(_04820_),
    .A3(_06867_),
    .B1(_06869_),
    .C1(_03459_),
    .Y(_06870_));
 sky130_fd_sc_hd__nor3_1 _25511_ (.A(_03460_),
    .B(_04852_),
    .C(_04863_),
    .Y(_06871_));
 sky130_fd_sc_hd__a211oi_1 _25512_ (.A1(_03460_),
    .A2(_04863_),
    .B1(_06871_),
    .C1(net3629),
    .Y(_06872_));
 sky130_fd_sc_hd__o22ai_2 _25513_ (.A1(_03800_),
    .A2(_06868_),
    .B1(_06870_),
    .B2(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__a21oi_1 _25514_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(_10746_),
    .B1(_03471_),
    .Y(_06874_));
 sky130_fd_sc_hd__nand3_1 _25515_ (.A(_10422_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .C(_03463_),
    .Y(_06875_));
 sky130_fd_sc_hd__o31ai_1 _25516_ (.A1(_10422_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A3(_03461_),
    .B1(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__a21oi_1 _25517_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(_03681_),
    .B1(_03463_),
    .Y(_06877_));
 sky130_fd_sc_hd__a21oi_1 _25518_ (.A1(_03681_),
    .A2(_06876_),
    .B1(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__o22ai_2 _25519_ (.A1(_03697_),
    .A2(_06874_),
    .B1(_06878_),
    .B2(_03471_),
    .Y(_06879_));
 sky130_fd_sc_hd__xnor2_1 _25520_ (.A(_03691_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__nor2_1 _25521_ (.A(_04051_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__and2_0 _25522_ (.A(_04051_),
    .B(_06880_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_1 _25523_ (.A(_06881_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__xnor2_1 _25524_ (.A(_06873_),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__xnor2_1 _25525_ (.A(_04608_),
    .B(_04873_),
    .Y(_06885_));
 sky130_fd_sc_hd__o221ai_1 _25526_ (.A1(_04651_),
    .A2(_04824_),
    .B1(_04873_),
    .B2(net3570),
    .C1(net3571),
    .Y(_06886_));
 sky130_fd_sc_hd__a221o_1 _25527_ (.A1(_04739_),
    .A2(_04824_),
    .B1(_04873_),
    .B2(_03951_),
    .C1(net3571),
    .X(_06887_));
 sky130_fd_sc_hd__nand3_1 _25528_ (.A(net3571),
    .B(_04828_),
    .C(_04873_),
    .Y(_06888_));
 sky130_fd_sc_hd__or3_1 _25529_ (.A(net3571),
    .B(_04828_),
    .C(_04873_),
    .X(_06889_));
 sky130_fd_sc_hd__a31oi_1 _25530_ (.A1(net3570),
    .A2(_06888_),
    .A3(_06889_),
    .B1(_04740_),
    .Y(_06890_));
 sky130_fd_sc_hd__a21oi_1 _25531_ (.A1(_06886_),
    .A2(_06887_),
    .B1(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2b_1 _25532_ (.A_N(_06891_),
    .B(_04859_),
    .Y(_06892_));
 sky130_fd_sc_hd__a21boi_4 _25533_ (.A1(_04739_),
    .A2(_06885_),
    .B1_N(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__xnor2_1 _25534_ (.A(_06884_),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__nor2_1 _25535_ (.A(_04839_),
    .B(_04842_),
    .Y(_06895_));
 sky130_fd_sc_hd__nand3_1 _25536_ (.A(net3632),
    .B(_02856_),
    .C(_04621_),
    .Y(_06896_));
 sky130_fd_sc_hd__o21ai_0 _25537_ (.A1(_02856_),
    .A2(_04621_),
    .B1(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__a21oi_1 _25538_ (.A1(_04621_),
    .A2(_04838_),
    .B1(net3632),
    .Y(_06898_));
 sky130_fd_sc_hd__nor3_1 _25539_ (.A(_02987_),
    .B(_06897_),
    .C(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__a21oi_1 _25540_ (.A1(_02987_),
    .A2(_03181_),
    .B1(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_1 _25541_ (.A(_04839_),
    .B(_04842_),
    .Y(_06901_));
 sky130_fd_sc_hd__a22oi_1 _25542_ (.A1(_04836_),
    .A2(_06901_),
    .B1(_06895_),
    .B2(_04621_),
    .Y(_06902_));
 sky130_fd_sc_hd__o221a_4 _25543_ (.A1(_04621_),
    .A2(_06895_),
    .B1(_06900_),
    .B2(_06902_),
    .C1(_04747_),
    .X(_06903_));
 sky130_fd_sc_hd__or2_4 _25544_ (.A(_06862_),
    .B(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__xnor2_1 _25545_ (.A(_04038_),
    .B(_04873_),
    .Y(_06905_));
 sky130_fd_sc_hd__nor2_1 _25546_ (.A(_03460_),
    .B(_04781_),
    .Y(_06906_));
 sky130_fd_sc_hd__nor2_1 _25547_ (.A(net3627),
    .B(_04855_),
    .Y(_06907_));
 sky130_fd_sc_hd__o21ai_0 _25548_ (.A1(_06906_),
    .A2(_06907_),
    .B1(net3629),
    .Y(_06908_));
 sky130_fd_sc_hd__o21ai_0 _25549_ (.A1(_03470_),
    .A2(_04855_),
    .B1(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__o21ai_0 _25550_ (.A1(net3627),
    .A2(_04781_),
    .B1(net3629),
    .Y(_06910_));
 sky130_fd_sc_hd__o21ai_0 _25551_ (.A1(_03460_),
    .A2(_04852_),
    .B1(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__nor3_1 _25552_ (.A(_04820_),
    .B(_04854_),
    .C(_06867_),
    .Y(_06912_));
 sky130_fd_sc_hd__a21oi_1 _25553_ (.A1(_06867_),
    .A2(_06911_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__nor2_1 _25554_ (.A(net3577),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__a31oi_2 _25555_ (.A1(net3577),
    .A2(_04863_),
    .A3(_06909_),
    .B1(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__o21ai_2 _25556_ (.A1(_03951_),
    .A2(_06905_),
    .B1(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__xnor2_1 _25557_ (.A(_04651_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__xnor2_1 _25558_ (.A(_06904_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__xnor2_2 _25559_ (.A(_06894_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__xor2_1 _25560_ (.A(_06866_),
    .B(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__xnor2_1 _25561_ (.A(_06863_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xnor2_1 _25562_ (.A(_06860_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__xnor2_1 _25563_ (.A(_06859_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__a21oi_1 _25564_ (.A1(_02000_),
    .A2(_06923_),
    .B1(_10690_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand2_1 _25565_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B(_06503_),
    .Y(_06925_));
 sky130_fd_sc_hd__o31ai_1 _25566_ (.A1(_06503_),
    .A2(_06852_),
    .A3(_06924_),
    .B1(_06925_),
    .Y(_01573_));
 sky130_fd_sc_hd__a31oi_1 _25567_ (.A1(_04345_),
    .A2(net3452),
    .A3(_04441_),
    .B1(_04381_),
    .Y(_06926_));
 sky130_fd_sc_hd__a21oi_1 _25568_ (.A1(_04345_),
    .A2(net3452),
    .B1(_04441_),
    .Y(_06927_));
 sky130_fd_sc_hd__clkinv_1 _25569_ (.A(_04885_),
    .Y(_06928_));
 sky130_fd_sc_hd__o211ai_1 _25570_ (.A1(_06926_),
    .A2(_06927_),
    .B1(_04562_),
    .C1(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2_1 _25571_ (.A(_04725_),
    .B(_06928_),
    .Y(_06930_));
 sky130_fd_sc_hd__xor2_1 _25572_ (.A(_06863_),
    .B(_06920_),
    .X(_06931_));
 sky130_fd_sc_hd__nand2_1 _25573_ (.A(_04809_),
    .B(_06853_),
    .Y(_06932_));
 sky130_fd_sc_hd__nor2_1 _25574_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__inv_1 _25575_ (.A(_06858_),
    .Y(_06934_));
 sky130_fd_sc_hd__o21ai_0 _25576_ (.A1(_06934_),
    .A2(_06931_),
    .B1(_06860_),
    .Y(_06935_));
 sky130_fd_sc_hd__a21boi_0 _25577_ (.A1(_04097_),
    .A2(net3458),
    .B1_N(_04251_),
    .Y(_06936_));
 sky130_fd_sc_hd__nand2_1 _25578_ (.A(_04254_),
    .B(_04345_),
    .Y(_06937_));
 sky130_fd_sc_hd__o2111ai_1 _25579_ (.A1(_06936_),
    .A2(_06937_),
    .B1(_04344_),
    .C1(_04597_),
    .D1(_06928_),
    .Y(_06938_));
 sky130_fd_sc_hd__nor2_1 _25580_ (.A(_04598_),
    .B(_04725_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_1 _25581_ (.A(_04885_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nor2_1 _25582_ (.A(_06932_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__a211o_1 _25583_ (.A1(_06938_),
    .A2(_06941_),
    .B1(_06858_),
    .C1(_06921_),
    .X(_06942_));
 sky130_fd_sc_hd__a32oi_2 _25584_ (.A1(_06929_),
    .A2(_06930_),
    .A3(_06933_),
    .B1(_06935_),
    .B2(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2b_1 _25585_ (.A_N(_06884_),
    .B(_06893_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2b_1 _25586_ (.A_N(_06893_),
    .B(_06884_),
    .Y(_06945_));
 sky130_fd_sc_hd__or3_1 _25587_ (.A(_04739_),
    .B(_06916_),
    .C(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__o21ai_0 _25588_ (.A1(_04651_),
    .A2(_06944_),
    .B1(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2b_1 _25589_ (.A_N(_06916_),
    .B(_06904_),
    .Y(_06948_));
 sky130_fd_sc_hd__nand2_1 _25590_ (.A(_04739_),
    .B(_06894_),
    .Y(_06949_));
 sky130_fd_sc_hd__o21ai_0 _25591_ (.A1(_04739_),
    .A2(_06944_),
    .B1(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__nor2_1 _25592_ (.A(_06884_),
    .B(_06916_),
    .Y(_06951_));
 sky130_fd_sc_hd__nor3b_1 _25593_ (.A(_06893_),
    .B(_06904_),
    .C_N(_06916_),
    .Y(_06952_));
 sky130_fd_sc_hd__a21oi_1 _25594_ (.A1(_06893_),
    .A2(_06951_),
    .B1(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__nand4b_1 _25595_ (.A_N(_06904_),
    .B(_06916_),
    .C(_06945_),
    .D(_04651_),
    .Y(_06954_));
 sky130_fd_sc_hd__o21ai_0 _25596_ (.A1(_04651_),
    .A2(_06953_),
    .B1(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__a221oi_1 _25597_ (.A1(_06904_),
    .A2(_06947_),
    .B1(_06948_),
    .B2(_06950_),
    .C1(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__a21oi_1 _25598_ (.A1(net3627),
    .A2(_04863_),
    .B1(net3629),
    .Y(_06957_));
 sky130_fd_sc_hd__a21oi_1 _25599_ (.A1(_03460_),
    .A2(_06867_),
    .B1(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand2_1 _25600_ (.A(_03803_),
    .B(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__a21oi_1 _25601_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A2(net3668),
    .B1(net3732),
    .Y(_06960_));
 sky130_fd_sc_hd__nand2_1 _25602_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B(net3668),
    .Y(_06961_));
 sky130_fd_sc_hd__nor2_1 _25603_ (.A(_03803_),
    .B(_06958_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand2b_1 _25604_ (.A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .Y(_06963_));
 sky130_fd_sc_hd__nand3b_1 _25605_ (.A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B(_06959_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_0 _25606_ (.A1(_06962_),
    .A2(_06963_),
    .B1(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__a22oi_1 _25607_ (.A1(_06961_),
    .A2(_06962_),
    .B1(_06965_),
    .B2(net3668),
    .Y(_06966_));
 sky130_fd_sc_hd__o22ai_1 _25608_ (.A1(_06959_),
    .A2(_06960_),
    .B1(_06966_),
    .B2(net3732),
    .Y(_06967_));
 sky130_fd_sc_hd__xnor2_1 _25609_ (.A(_06903_),
    .B(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__nor3_1 _25610_ (.A(_04051_),
    .B(_06873_),
    .C(_06880_),
    .Y(_06969_));
 sky130_fd_sc_hd__a21oi_1 _25611_ (.A1(_06873_),
    .A2(_06882_),
    .B1(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__xnor2_1 _25612_ (.A(_06968_),
    .B(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__xnor2_1 _25613_ (.A(_06956_),
    .B(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand2_1 _25614_ (.A(_06863_),
    .B(_06919_),
    .Y(_06973_));
 sky130_fd_sc_hd__nor2_1 _25615_ (.A(_06863_),
    .B(_06919_),
    .Y(_06974_));
 sky130_fd_sc_hd__a21oi_2 _25616_ (.A1(_06866_),
    .A2(_06973_),
    .B1(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__xnor2_1 _25617_ (.A(_06972_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__xnor2_1 _25618_ (.A(_06943_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__nor2b_1 _25619_ (.A(_06503_),
    .B_N(_06851_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_0 _25620_ (.A1(_10690_),
    .A2(_06977_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__nand2_1 _25621_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B(_06503_),
    .Y(_06980_));
 sky130_fd_sc_hd__nand2_1 _25622_ (.A(_06979_),
    .B(_06980_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _25623_ (.A(net3529),
    .B(_02990_),
    .Y(_06981_));
 sky130_fd_sc_hd__a21oi_1 _25624_ (.A1(net3727),
    .A2(_02990_),
    .B1(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_1 _25625_ (.A(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .B(_06384_),
    .Y(_06983_));
 sky130_fd_sc_hd__o21ai_0 _25626_ (.A1(_10684_),
    .A2(_06982_),
    .B1(_06983_),
    .Y(_01575_));
 sky130_fd_sc_hd__mux2i_1 _25627_ (.A0(net3530),
    .A1(_08777_),
    .S(_04421_),
    .Y(_06984_));
 sky130_fd_sc_hd__nand2_1 _25628_ (.A(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .B(_06384_),
    .Y(_06985_));
 sky130_fd_sc_hd__o21ai_0 _25629_ (.A1(_10684_),
    .A2(_06984_),
    .B1(_06985_),
    .Y(_01576_));
 sky130_fd_sc_hd__mux2i_1 _25630_ (.A0(net3519),
    .A1(_08917_),
    .S(_04421_),
    .Y(_06986_));
 sky130_fd_sc_hd__nand2_1 _25631_ (.A(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .B(_06384_),
    .Y(_06987_));
 sky130_fd_sc_hd__o21ai_0 _25632_ (.A1(_10684_),
    .A2(_06986_),
    .B1(_06987_),
    .Y(_01577_));
 sky130_fd_sc_hd__mux2i_1 _25633_ (.A0(net3520),
    .A1(net3706),
    .S(_04421_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_1 _25634_ (.A(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .B(_06384_),
    .Y(_06989_));
 sky130_fd_sc_hd__o21ai_0 _25635_ (.A1(_10684_),
    .A2(_06988_),
    .B1(_06989_),
    .Y(_01578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_83 ();
 sky130_fd_sc_hd__nor2b_4 _25637_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B_N(net59),
    .Y(_06991_));
 sky130_fd_sc_hd__nand2_2 _25638_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(_07869_),
    .Y(_06992_));
 sky130_fd_sc_hd__nor2_2 _25639_ (.A(net25),
    .B(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__nand2_1 _25640_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .B(net59),
    .Y(_06994_));
 sky130_fd_sc_hd__nor2_1 _25641_ (.A(net25),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__a31oi_1 _25642_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(\load_store_unit_i.ls_fsm_cs[1] ),
    .A3(\load_store_unit_i.lsu_err_q ),
    .B1(\load_store_unit_i.ls_fsm_cs[2] ),
    .Y(_06996_));
 sky130_fd_sc_hd__o21ai_0 _25643_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_06995_),
    .B1(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__a21boi_2 _25644_ (.A1(_10659_),
    .A2(_06997_),
    .B1_N(net26),
    .Y(_06998_));
 sky130_fd_sc_hd__a21oi_4 _25645_ (.A1(_06991_),
    .A2(_06993_),
    .B1(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_81 ();
 sky130_fd_sc_hd__nand2_1 _25648_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .B(_06999_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21ai_0 _25649_ (.A1(_10701_),
    .A2(_06999_),
    .B1(_07002_),
    .Y(_01580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_80 ();
 sky130_fd_sc_hd__mux2_1 _25651_ (.A0(net3515),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .S(net3555),
    .X(_01581_));
 sky130_fd_sc_hd__nor2_1 _25652_ (.A(net152),
    .B(net3555),
    .Y(_07004_));
 sky130_fd_sc_hd__a21oi_1 _25653_ (.A1(_08986_),
    .A2(net3555),
    .B1(_07004_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_4 _25654_ (.A(net3514),
    .B(_06999_),
    .Y(_07005_));
 sky130_fd_sc_hd__a21oi_1 _25655_ (.A1(_09212_),
    .A2(net3555),
    .B1(_07005_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _25656_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .B(net3555),
    .Y(_07006_));
 sky130_fd_sc_hd__o21ai_0 _25657_ (.A1(net3498),
    .A2(net3555),
    .B1(_07006_),
    .Y(_01584_));
 sky130_fd_sc_hd__mux2_1 _25658_ (.A0(net3513),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .S(net3555),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _25659_ (.A0(net3507),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .S(net3555),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _25660_ (.A0(net3506),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .S(net3555),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _25661_ (.A0(net3512),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .S(net3555),
    .X(_01588_));
 sky130_fd_sc_hd__inv_1 _25662_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .Y(_07007_));
 sky130_fd_sc_hd__mux2i_1 _25663_ (.A0(net3497),
    .A1(_07007_),
    .S(net3555),
    .Y(_01589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_79 ();
 sky130_fd_sc_hd__mux2_1 _25665_ (.A0(net160),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .S(net3555),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _25666_ (.A0(_06418_),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .S(net3555),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _25667_ (.A0(net161),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .S(net3555),
    .X(_01592_));
 sky130_fd_sc_hd__nand2_1 _25668_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .B(net3555),
    .Y(_07009_));
 sky130_fd_sc_hd__o21ai_0 _25669_ (.A1(net3496),
    .A2(net3555),
    .B1(_07009_),
    .Y(_01593_));
 sky130_fd_sc_hd__mux2_1 _25670_ (.A0(net3503),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .S(net3555),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _25671_ (.A0(net164),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .S(net3555),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _25672_ (.A0(net273),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .S(net3555),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _25673_ (.A0(net3495),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .S(net3555),
    .X(_01597_));
 sky130_fd_sc_hd__nand2_1 _25674_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .B(net3555),
    .Y(_07010_));
 sky130_fd_sc_hd__o21ai_0 _25675_ (.A1(net3486),
    .A2(net3555),
    .B1(_07010_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _25676_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .B(net3555),
    .Y(_07011_));
 sky130_fd_sc_hd__o21ai_0 _25677_ (.A1(net3487),
    .A2(net3555),
    .B1(_07011_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_1 _25678_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .B(net3555),
    .Y(_07012_));
 sky130_fd_sc_hd__o21ai_0 _25679_ (.A1(net3485),
    .A2(net3555),
    .B1(_07012_),
    .Y(_01600_));
 sky130_fd_sc_hd__mux2_1 _25680_ (.A0(net3474),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .S(net3555),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _25681_ (.A0(net3549),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .S(_06999_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _25682_ (.A0(net3473),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .S(net3555),
    .X(_01603_));
 sky130_fd_sc_hd__nand2_1 _25683_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .B(net3555),
    .Y(_07013_));
 sky130_fd_sc_hd__o21ai_0 _25684_ (.A1(net3471),
    .A2(net3555),
    .B1(_07013_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _25685_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .B(net3555),
    .Y(_07014_));
 sky130_fd_sc_hd__o21ai_0 _25686_ (.A1(net3534),
    .A2(net3555),
    .B1(_07014_),
    .Y(_01605_));
 sky130_fd_sc_hd__mux2_1 _25687_ (.A0(net3535),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .S(_06999_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _25688_ (.A0(net3537),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .S(net3555),
    .X(_01607_));
 sky130_fd_sc_hd__nand2_1 _25689_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .B(_06999_),
    .Y(_07015_));
 sky130_fd_sc_hd__o21ai_0 _25690_ (.A1(net3529),
    .A2(_06999_),
    .B1(_07015_),
    .Y(_01608_));
 sky130_fd_sc_hd__mux2_1 _25691_ (.A0(net3530),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .S(net3555),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _25692_ (.A0(net3519),
    .A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .S(_06999_),
    .X(_01610_));
 sky130_fd_sc_hd__nor2_1 _25693_ (.A(net3520),
    .B(net3555),
    .Y(_07016_));
 sky130_fd_sc_hd__a21oi_1 _25694_ (.A1(_08888_),
    .A2(net3555),
    .B1(_07016_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2b_1 _25695_ (.A(_10662_),
    .B_N(\load_store_unit_i.data_sign_ext_q ),
    .Y(_07017_));
 sky130_fd_sc_hd__a41o_1 _25696_ (.A1(_08009_),
    .A2(_07883_),
    .A3(_08005_),
    .A4(_10662_),
    .B1(_07017_),
    .X(_01612_));
 sky130_fd_sc_hd__and3_4 _25697_ (.A(net3831),
    .B(net3753),
    .C(_10536_),
    .X(net218));
 sky130_fd_sc_hd__nand2_1 _25698_ (.A(_10662_),
    .B(net218),
    .Y(_07018_));
 sky130_fd_sc_hd__o21ai_0 _25699_ (.A1(_10651_),
    .A2(_10662_),
    .B1(_07018_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _25700_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_07019_));
 sky130_fd_sc_hd__nand2_1 _25701_ (.A(_10657_),
    .B(_10658_),
    .Y(_07020_));
 sky130_fd_sc_hd__nand2_1 _25702_ (.A(_07019_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__nand2_2 _25703_ (.A(_10660_),
    .B(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__a21oi_1 _25704_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_06991_),
    .B1(net26),
    .Y(_07023_));
 sky130_fd_sc_hd__nand2b_4 _25705_ (.A_N(net3938),
    .B(net3753),
    .Y(_07024_));
 sky130_fd_sc_hd__a21oi_1 _25706_ (.A1(net3941),
    .A2(_06418_),
    .B1(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__nor2_1 _25707_ (.A(_10701_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__a21oi_2 _25708_ (.A1(_07024_),
    .A2(_06418_),
    .B1(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__o21ai_0 _25709_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_07019_),
    .B1(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand3_1 _25710_ (.A(_10660_),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .C(net26),
    .Y(_07029_));
 sky130_fd_sc_hd__nand2_1 _25711_ (.A(_07028_),
    .B(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__o21ai_0 _25712_ (.A1(_07022_),
    .A2(_07023_),
    .B1(\load_store_unit_i.handle_misaligned_q ),
    .Y(_07031_));
 sky130_fd_sc_hd__o31ai_1 _25713_ (.A1(_07022_),
    .A2(_07023_),
    .A3(_07030_),
    .B1(_07031_),
    .Y(_01614_));
 sky130_fd_sc_hd__o21ai_0 _25714_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_07020_),
    .B1(_06994_),
    .Y(_07032_));
 sky130_fd_sc_hd__nor2_1 _25715_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nor3_1 _25716_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(net26),
    .C(_07033_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2b_1 _25717_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B_N(_07027_),
    .Y(_07034_));
 sky130_fd_sc_hd__inv_1 _25718_ (.A(_07022_),
    .Y(net185));
 sky130_fd_sc_hd__o21ai_0 _25719_ (.A1(net26),
    .A2(_07034_),
    .B1(net185),
    .Y(_07035_));
 sky130_fd_sc_hd__a22oi_1 _25720_ (.A1(net59),
    .A2(_07022_),
    .B1(_07027_),
    .B2(net26),
    .Y(_07036_));
 sky130_fd_sc_hd__a21oi_1 _25721_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(net26),
    .B1(\load_store_unit_i.ls_fsm_cs[2] ),
    .Y(_07037_));
 sky130_fd_sc_hd__o21ai_0 _25722_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_07036_),
    .B1(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21oi_1 _25723_ (.A1(_07869_),
    .A2(_07035_),
    .B1(_07038_),
    .Y(_01616_));
 sky130_fd_sc_hd__a211oi_1 _25724_ (.A1(_06992_),
    .A2(_07029_),
    .B1(\load_store_unit_i.ls_fsm_cs[0] ),
    .C1(net59),
    .Y(_01617_));
 sky130_fd_sc_hd__inv_1 _25725_ (.A(net25),
    .Y(_07039_));
 sky130_fd_sc_hd__xor2_1 _25726_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .X(_07040_));
 sky130_fd_sc_hd__nand2_2 _25727_ (.A(_06991_),
    .B(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__nand3_1 _25728_ (.A(\load_store_unit_i.lsu_err_q ),
    .B(_10659_),
    .C(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__o21ai_0 _25729_ (.A1(_07039_),
    .A2(_07041_),
    .B1(_07042_),
    .Y(_01618_));
 sky130_fd_sc_hd__mux2i_1 _25730_ (.A0(_02419_),
    .A1(_10701_),
    .S(_10662_),
    .Y(_01619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_78 ();
 sky130_fd_sc_hd__nor2_1 _25732_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_10662_),
    .Y(_07044_));
 sky130_fd_sc_hd__a21oi_1 _25733_ (.A1(_10662_),
    .A2(net3562),
    .B1(_07044_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_4 _25734_ (.A(\load_store_unit_i.data_we_q ),
    .B(_07041_),
    .Y(_07045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__mux2_1 _25736_ (.A0(\load_store_unit_i.rdata_q[0] ),
    .A1(net57),
    .S(net3729),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _25737_ (.A0(\load_store_unit_i.rdata_q[10] ),
    .A1(net36),
    .S(net3729),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _25738_ (.A0(\load_store_unit_i.rdata_q[11] ),
    .A1(net37),
    .S(_07045_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _25739_ (.A0(\load_store_unit_i.rdata_q[12] ),
    .A1(net39),
    .S(_07045_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _25740_ (.A0(\load_store_unit_i.rdata_q[13] ),
    .A1(net40),
    .S(net3729),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _25741_ (.A0(\load_store_unit_i.rdata_q[14] ),
    .A1(net41),
    .S(_07045_),
    .X(_01626_));
 sky130_fd_sc_hd__nand2_1 _25742_ (.A(net42),
    .B(_07045_),
    .Y(_07047_));
 sky130_fd_sc_hd__o21ai_0 _25743_ (.A1(_02845_),
    .A2(_07045_),
    .B1(_07047_),
    .Y(_01627_));
 sky130_fd_sc_hd__mux2_1 _25744_ (.A0(\load_store_unit_i.rdata_q[16] ),
    .A1(net43),
    .S(net3729),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _25745_ (.A0(\load_store_unit_i.rdata_q[17] ),
    .A1(net44),
    .S(net3729),
    .X(_01629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__mux2_1 _25747_ (.A0(\load_store_unit_i.rdata_q[18] ),
    .A1(net45),
    .S(net3729),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _25748_ (.A0(\load_store_unit_i.rdata_q[19] ),
    .A1(net46),
    .S(net3729),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _25749_ (.A0(\load_store_unit_i.rdata_q[1] ),
    .A1(net58),
    .S(net3729),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _25750_ (.A0(\load_store_unit_i.rdata_q[20] ),
    .A1(net47),
    .S(_07045_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _25751_ (.A0(\load_store_unit_i.rdata_q[21] ),
    .A1(net48),
    .S(_07045_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _25752_ (.A0(\load_store_unit_i.rdata_q[22] ),
    .A1(net50),
    .S(_07045_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _25753_ (.A0(\load_store_unit_i.rdata_q[23] ),
    .A1(net51),
    .S(_07045_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _25754_ (.A0(\load_store_unit_i.rdata_q[2] ),
    .A1(net28),
    .S(net3729),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _25755_ (.A0(\load_store_unit_i.rdata_q[3] ),
    .A1(net29),
    .S(_07045_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _25756_ (.A0(\load_store_unit_i.rdata_q[4] ),
    .A1(net30),
    .S(_07045_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _25757_ (.A0(\load_store_unit_i.rdata_q[5] ),
    .A1(net31),
    .S(net3729),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _25758_ (.A0(\load_store_unit_i.rdata_q[6] ),
    .A1(net32),
    .S(_07045_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _25759_ (.A0(\load_store_unit_i.rdata_q[7] ),
    .A1(net33),
    .S(_07045_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _25760_ (.A0(\load_store_unit_i.rdata_q[8] ),
    .A1(net34),
    .S(net3729),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _25761_ (.A0(\load_store_unit_i.rdata_q[9] ),
    .A1(net35),
    .S(_07045_),
    .X(_01644_));
 sky130_fd_sc_hd__inv_1 _25762_ (.A(_12393_),
    .Y(_07049_));
 sky130_fd_sc_hd__and2_4 _25763_ (.A(_10595_),
    .B(net3501),
    .X(_07050_));
 sky130_fd_sc_hd__nand3_1 _25764_ (.A(_11177_),
    .B(_11197_),
    .C(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__a22oi_1 _25765_ (.A1(net3545),
    .A2(_07049_),
    .B1(_12476_),
    .B2(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__nor2_1 _25766_ (.A(\cs_registers_i.mstatus_q[2] ),
    .B(_07050_),
    .Y(_07053_));
 sky130_fd_sc_hd__a22oi_1 _25767_ (.A1(net3950),
    .A2(net3532),
    .B1(_12400_),
    .B2(\cs_registers_i.mstack_q[0] ),
    .Y(_07054_));
 sky130_fd_sc_hd__o21ai_0 _25768_ (.A1(_07052_),
    .A2(_07053_),
    .B1(_07054_),
    .Y(_00383_));
 sky130_fd_sc_hd__nor2_1 _25769_ (.A(\cs_registers_i.mstatus_q[3] ),
    .B(_07050_),
    .Y(_07055_));
 sky130_fd_sc_hd__a22oi_1 _25770_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(_12394_),
    .B1(_12400_),
    .B2(\cs_registers_i.mstack_q[1] ),
    .Y(_07056_));
 sky130_fd_sc_hd__o21ai_0 _25771_ (.A1(_07052_),
    .A2(_07055_),
    .B1(_07056_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2b_1 _25772_ (.A_N(\cs_registers_i.mstack_q[2] ),
    .B(\cs_registers_i.nmi_mode_i ),
    .Y(_07057_));
 sky130_fd_sc_hd__and3_4 _25773_ (.A(_10541_),
    .B(_10545_),
    .C(_10586_),
    .X(_07058_));
 sky130_fd_sc_hd__nand4_1 _25774_ (.A(_11014_),
    .B(_10634_),
    .C(_10589_),
    .D(_07058_),
    .Y(_07059_));
 sky130_fd_sc_hd__a22o_1 _25775_ (.A1(net3545),
    .A2(_07049_),
    .B1(_12476_),
    .B2(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__a222oi_1 _25776_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(net3532),
    .B1(net3663),
    .B2(_07057_),
    .C1(_07060_),
    .C2(\cs_registers_i.mstatus_q[4] ),
    .Y(_07061_));
 sky130_fd_sc_hd__o21ai_0 _25777_ (.A1(_11685_),
    .A2(_12744_),
    .B1(_07061_),
    .Y(_00385_));
 sky130_fd_sc_hd__a22oi_1 _25778_ (.A1(\cs_registers_i.mstatus_q[4] ),
    .A2(net3663),
    .B1(_07060_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .Y(_07062_));
 sky130_fd_sc_hd__o21ai_0 _25779_ (.A1(_11612_),
    .A2(_12744_),
    .B1(_07062_),
    .Y(_00386_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__nand2_1 _25781_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .Y(_07064_));
 sky130_fd_sc_hd__nand3_1 _25782_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_10908_),
    .C(net94),
    .Y(_07065_));
 sky130_fd_sc_hd__nand2b_1 _25783_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .B(net3948),
    .Y(_07066_));
 sky130_fd_sc_hd__a21oi_1 _25784_ (.A1(_07064_),
    .A2(_07065_),
    .B1(_07066_),
    .Y(_01579_));
 sky130_fd_sc_hd__o21ai_2 _25785_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B1(_10798_),
    .Y(_07067_));
 sky130_fd_sc_hd__o21ai_0 _25786_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_07068_));
 sky130_fd_sc_hd__nor2_2 _25787_ (.A(_10826_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__a211oi_4 _25788_ (.A1(_10538_),
    .A2(_07067_),
    .B1(_07069_),
    .C1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_07070_));
 sky130_fd_sc_hd__nor2_2 _25789_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__nor4b_1 _25790_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .B(_10978_),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .D_N(_10653_),
    .Y(_07072_));
 sky130_fd_sc_hd__o211ai_1 _25791_ (.A1(_10495_),
    .A2(_06350_),
    .B1(_07071_),
    .C1(_07072_),
    .Y(core_busy_d));
 sky130_fd_sc_hd__and2_1 _25792_ (.A(clknet_1_0__leaf_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .X(clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__nand2_1 _25794_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B(_07024_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand2_1 _25795_ (.A(net3753),
    .B(_10510_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand2_1 _25796_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__a21oi_1 _25797_ (.A1(_10701_),
    .A2(net3562),
    .B1(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__a31o_1 _25798_ (.A1(_10701_),
    .A2(net3562),
    .A3(_07074_),
    .B1(_07077_),
    .X(net181));
 sky130_fd_sc_hd__nand3_1 _25799_ (.A(net3753),
    .B(_10510_),
    .C(_10701_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand3_1 _25800_ (.A(net3562),
    .B(_07076_),
    .C(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__o21ai_0 _25801_ (.A1(net3562),
    .A2(_07074_),
    .B1(_07079_),
    .Y(net182));
 sky130_fd_sc_hd__nor2_1 _25802_ (.A(_08008_),
    .B(_10701_),
    .Y(_07080_));
 sky130_fd_sc_hd__o21ai_0 _25803_ (.A1(_07024_),
    .A2(_07080_),
    .B1(net3562),
    .Y(_07081_));
 sky130_fd_sc_hd__nor2_1 _25804_ (.A(_10701_),
    .B(_07074_),
    .Y(_07082_));
 sky130_fd_sc_hd__a21oi_1 _25805_ (.A1(_10701_),
    .A2(_07076_),
    .B1(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__o22ai_1 _25806_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_07081_),
    .B1(_07083_),
    .B2(net3562),
    .Y(net183));
 sky130_fd_sc_hd__o32ai_1 _25807_ (.A1(_07075_),
    .A2(_10701_),
    .A3(net3562),
    .B1(_07025_),
    .B2(\load_store_unit_i.handle_misaligned_q ),
    .Y(net184));
 sky130_fd_sc_hd__mux2i_1 _25808_ (.A0(_08917_),
    .A1(_10010_),
    .S(net3562),
    .Y(_07084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__nand2_1 _25810_ (.A(net3712),
    .B(net3562),
    .Y(_07086_));
 sky130_fd_sc_hd__o21ai_0 _25811_ (.A1(_09489_),
    .A2(net3562),
    .B1(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__mux2i_1 _25812_ (.A0(_07084_),
    .A1(_07087_),
    .S(net3575),
    .Y(net186));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__mux2i_1 _25814_ (.A0(net3715),
    .A1(net3692),
    .S(net3556),
    .Y(_07089_));
 sky130_fd_sc_hd__mux2i_1 _25815_ (.A0(net3701),
    .A1(net3683),
    .S(net3556),
    .Y(_07090_));
 sky130_fd_sc_hd__mux2i_1 _25816_ (.A0(_07089_),
    .A1(_07090_),
    .S(net3575),
    .Y(net187));
 sky130_fd_sc_hd__mux2i_1 _25817_ (.A0(net3719),
    .A1(_09564_),
    .S(net3556),
    .Y(_07091_));
 sky130_fd_sc_hd__nand2_1 _25818_ (.A(net3680),
    .B(net3556),
    .Y(_07092_));
 sky130_fd_sc_hd__o21ai_0 _25819_ (.A1(net261),
    .A2(net3556),
    .B1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__mux2i_1 _25820_ (.A0(_07091_),
    .A1(_07093_),
    .S(net3575),
    .Y(net188));
 sky130_fd_sc_hd__mux2i_1 _25821_ (.A0(net3707),
    .A1(net3688),
    .S(net3556),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_1 _25822_ (.A(_09243_),
    .B(net3562),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_1 _25823_ (.A(_10294_),
    .B(net3556),
    .Y(_07096_));
 sky130_fd_sc_hd__nand2_1 _25824_ (.A(_07095_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__mux2i_1 _25825_ (.A0(_07094_),
    .A1(_07097_),
    .S(net3575),
    .Y(net189));
 sky130_fd_sc_hd__mux2i_1 _25826_ (.A0(_08240_),
    .A1(net3691),
    .S(net3556),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_1 _25827_ (.A(_09149_),
    .B(net3562),
    .Y(_07099_));
 sky130_fd_sc_hd__o21ai_0 _25828_ (.A1(_10360_),
    .A2(net3562),
    .B1(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__mux2i_1 _25829_ (.A0(_07098_),
    .A1(_07100_),
    .S(net3575),
    .Y(net190));
 sky130_fd_sc_hd__mux2i_1 _25830_ (.A0(net3727),
    .A1(net3686),
    .S(net3556),
    .Y(_07101_));
 sky130_fd_sc_hd__mux2i_1 _25831_ (.A0(net3696),
    .A1(_10474_),
    .S(net3556),
    .Y(_07102_));
 sky130_fd_sc_hd__mux2i_1 _25832_ (.A0(_07101_),
    .A1(_07102_),
    .S(net3575),
    .Y(net191));
 sky130_fd_sc_hd__mux2i_1 _25833_ (.A0(net425),
    .A1(net3685),
    .S(net3556),
    .Y(_07103_));
 sky130_fd_sc_hd__o21a_4 _25834_ (.A1(net3849),
    .A2(_09267_),
    .B1(_09275_),
    .X(_07104_));
 sky130_fd_sc_hd__nand2_1 _25835_ (.A(_10390_),
    .B(net3556),
    .Y(_07105_));
 sky130_fd_sc_hd__o21ai_0 _25836_ (.A1(_07104_),
    .A2(net3556),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__mux2i_1 _25837_ (.A0(_07103_),
    .A1(_07106_),
    .S(net3575),
    .Y(net192));
 sky130_fd_sc_hd__mux2i_1 _25838_ (.A0(_08917_),
    .A1(_10010_),
    .S(net3556),
    .Y(_07107_));
 sky130_fd_sc_hd__nand2_1 _25839_ (.A(net3712),
    .B(net3556),
    .Y(_07108_));
 sky130_fd_sc_hd__o21ai_0 _25840_ (.A1(_09489_),
    .A2(net3556),
    .B1(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__mux2i_1 _25841_ (.A0(_07107_),
    .A1(_07109_),
    .S(net3575),
    .Y(net193));
 sky130_fd_sc_hd__nand2_1 _25842_ (.A(_10062_),
    .B(net3556),
    .Y(_07110_));
 sky130_fd_sc_hd__o21ai_0 _25843_ (.A1(net3706),
    .A2(net3556),
    .B1(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand2_1 _25844_ (.A(net342),
    .B(net3556),
    .Y(_07112_));
 sky130_fd_sc_hd__o21ai_0 _25845_ (.A1(net409),
    .A2(net3556),
    .B1(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__mux2i_1 _25847_ (.A0(_07111_),
    .A1(_07113_),
    .S(net3575),
    .Y(net194));
 sky130_fd_sc_hd__mux2i_1 _25848_ (.A0(net3715),
    .A1(net3692),
    .S(net3562),
    .Y(_07115_));
 sky130_fd_sc_hd__mux2i_1 _25849_ (.A0(_07090_),
    .A1(_07115_),
    .S(net3575),
    .Y(net195));
 sky130_fd_sc_hd__mux2i_1 _25850_ (.A0(net3719),
    .A1(_09564_),
    .S(net3562),
    .Y(_07116_));
 sky130_fd_sc_hd__mux2i_1 _25851_ (.A0(_07093_),
    .A1(_07116_),
    .S(net3575),
    .Y(net196));
 sky130_fd_sc_hd__nor2_1 _25852_ (.A(_10062_),
    .B(net3556),
    .Y(_07117_));
 sky130_fd_sc_hd__a21oi_1 _25853_ (.A1(net3706),
    .A2(net3556),
    .B1(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__nand2_1 _25854_ (.A(net342),
    .B(net3562),
    .Y(_07119_));
 sky130_fd_sc_hd__o21ai_0 _25855_ (.A1(net409),
    .A2(net3562),
    .B1(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__mux2i_1 _25856_ (.A0(_07118_),
    .A1(_07120_),
    .S(net3575),
    .Y(net197));
 sky130_fd_sc_hd__mux2i_1 _25857_ (.A0(net3707),
    .A1(net3688),
    .S(net3562),
    .Y(_07121_));
 sky130_fd_sc_hd__mux2i_1 _25858_ (.A0(_07097_),
    .A1(_07121_),
    .S(net3575),
    .Y(net198));
 sky130_fd_sc_hd__mux2i_1 _25859_ (.A0(_08240_),
    .A1(net3691),
    .S(net3562),
    .Y(_07122_));
 sky130_fd_sc_hd__mux2i_1 _25860_ (.A0(_07100_),
    .A1(_07122_),
    .S(net3575),
    .Y(net199));
 sky130_fd_sc_hd__mux2i_1 _25861_ (.A0(net3727),
    .A1(net3686),
    .S(net3562),
    .Y(_07123_));
 sky130_fd_sc_hd__mux2i_1 _25862_ (.A0(_07102_),
    .A1(_07123_),
    .S(net3575),
    .Y(net200));
 sky130_fd_sc_hd__mux2i_1 _25863_ (.A0(net425),
    .A1(net3685),
    .S(net3562),
    .Y(_07124_));
 sky130_fd_sc_hd__mux2i_1 _25864_ (.A0(_07106_),
    .A1(_07124_),
    .S(net3575),
    .Y(net201));
 sky130_fd_sc_hd__mux2i_1 _25865_ (.A0(_07109_),
    .A1(_07084_),
    .S(net3575),
    .Y(net202));
 sky130_fd_sc_hd__mux2i_1 _25866_ (.A0(_07113_),
    .A1(_07118_),
    .S(net3575),
    .Y(net203));
 sky130_fd_sc_hd__mux2i_1 _25867_ (.A0(net3701),
    .A1(net3683),
    .S(net3562),
    .Y(_07125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__mux2i_1 _25869_ (.A0(_07115_),
    .A1(_07125_),
    .S(net3575),
    .Y(net204));
 sky130_fd_sc_hd__nand2_1 _25870_ (.A(net3680),
    .B(net3562),
    .Y(_07127_));
 sky130_fd_sc_hd__o21ai_0 _25871_ (.A1(net261),
    .A2(net3562),
    .B1(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__mux2i_1 _25872_ (.A0(_07116_),
    .A1(_07128_),
    .S(net3575),
    .Y(net205));
 sky130_fd_sc_hd__nand2_1 _25873_ (.A(_10294_),
    .B(net3562),
    .Y(_07129_));
 sky130_fd_sc_hd__nand2_1 _25874_ (.A(_09243_),
    .B(net3556),
    .Y(_07130_));
 sky130_fd_sc_hd__nand2_1 _25875_ (.A(_07129_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__mux2i_1 _25876_ (.A0(_07121_),
    .A1(_07131_),
    .S(net3575),
    .Y(net206));
 sky130_fd_sc_hd__nand2_1 _25877_ (.A(_09149_),
    .B(net3556),
    .Y(_07132_));
 sky130_fd_sc_hd__o21ai_0 _25878_ (.A1(_10360_),
    .A2(net3556),
    .B1(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__mux2i_1 _25879_ (.A0(_07122_),
    .A1(_07133_),
    .S(net3575),
    .Y(net207));
 sky130_fd_sc_hd__mux2i_1 _25880_ (.A0(_07125_),
    .A1(_07089_),
    .S(net3575),
    .Y(net208));
 sky130_fd_sc_hd__mux2i_1 _25881_ (.A0(net3696),
    .A1(_10474_),
    .S(net3562),
    .Y(_07134_));
 sky130_fd_sc_hd__mux2i_1 _25882_ (.A0(_07123_),
    .A1(_07134_),
    .S(net3575),
    .Y(net209));
 sky130_fd_sc_hd__nand2_1 _25883_ (.A(_10390_),
    .B(net3562),
    .Y(_07135_));
 sky130_fd_sc_hd__o21ai_0 _25884_ (.A1(_07104_),
    .A2(net3562),
    .B1(_07135_),
    .Y(_07136_));
 sky130_fd_sc_hd__mux2i_1 _25885_ (.A0(_07124_),
    .A1(_07136_),
    .S(net3575),
    .Y(net210));
 sky130_fd_sc_hd__mux2i_1 _25886_ (.A0(_07128_),
    .A1(_07091_),
    .S(net3575),
    .Y(net211));
 sky130_fd_sc_hd__mux2i_1 _25887_ (.A0(_07131_),
    .A1(_07094_),
    .S(net3575),
    .Y(net212));
 sky130_fd_sc_hd__mux2i_1 _25888_ (.A0(_07133_),
    .A1(_07098_),
    .S(net3575),
    .Y(net213));
 sky130_fd_sc_hd__mux2i_1 _25889_ (.A0(_07134_),
    .A1(_07101_),
    .S(net3575),
    .Y(net214));
 sky130_fd_sc_hd__mux2i_1 _25890_ (.A0(_07136_),
    .A1(_07103_),
    .S(net3575),
    .Y(net215));
 sky130_fd_sc_hd__mux2i_1 _25891_ (.A0(_07087_),
    .A1(_07107_),
    .S(net3575),
    .Y(net216));
 sky130_fd_sc_hd__mux2i_1 _25892_ (.A0(_07120_),
    .A1(_07111_),
    .S(net3575),
    .Y(net217));
 sky130_fd_sc_hd__nand2_8 _25893_ (.A(_10769_),
    .B(_10775_),
    .Y(_07137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_69 ();
 sky130_fd_sc_hd__nand2_1 _25895_ (.A(_10858_),
    .B(_10862_),
    .Y(_07139_));
 sky130_fd_sc_hd__nand2_8 _25896_ (.A(_10872_),
    .B(_10879_),
    .Y(_07140_));
 sky130_fd_sc_hd__nor2_4 _25897_ (.A(_10867_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_68 ();
 sky130_fd_sc_hd__nor3_2 _25899_ (.A(_10866_),
    .B(_10872_),
    .C(_10879_),
    .Y(_07143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__nand2_4 _25901_ (.A(_10838_),
    .B(_10842_),
    .Y(_07145_));
 sky130_fd_sc_hd__or4_4 _25902_ (.A(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .B(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .C(_10892_),
    .D(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__nor2_1 _25903_ (.A(_10898_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__a32oi_1 _25904_ (.A1(_10898_),
    .A2(_07139_),
    .A3(_07141_),
    .B1(_07143_),
    .B2(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_66 ();
 sky130_fd_sc_hd__nand2_8 _25906_ (.A(net3733),
    .B(_10873_),
    .Y(_07150_));
 sky130_fd_sc_hd__nor2_4 _25907_ (.A(_10769_),
    .B(_10776_),
    .Y(_07151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__nand2_1 _25909_ (.A(_07150_),
    .B(_07151_),
    .Y(_07153_));
 sky130_fd_sc_hd__nor4_2 _25910_ (.A(\if_stage_i.compressed_decoder_i.instr_i[7] ),
    .B(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .C(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .D(_10862_),
    .Y(_07154_));
 sky130_fd_sc_hd__nor2b_4 _25911_ (.A(_10850_),
    .B_N(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__nor2_2 _25912_ (.A(_10898_),
    .B(_07145_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_8 _25913_ (.A(_10866_),
    .B(_10878_),
    .Y(_07157_));
 sky130_fd_sc_hd__a21oi_1 _25914_ (.A1(_07155_),
    .A2(_07156_),
    .B1(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_4 _25915_ (.A(_10867_),
    .B(_10879_),
    .Y(_07159_));
 sky130_fd_sc_hd__nand2_8 _25916_ (.A(_10872_),
    .B(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_63 ();
 sky130_fd_sc_hd__nor2_4 _25919_ (.A(_10769_),
    .B(_10775_),
    .Y(_07163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_61 ();
 sky130_fd_sc_hd__a21oi_1 _25922_ (.A1(_07155_),
    .A2(_07147_),
    .B1(_10878_),
    .Y(_07166_));
 sky130_fd_sc_hd__a21oi_1 _25923_ (.A1(_10878_),
    .A2(_07155_),
    .B1(_10867_),
    .Y(_07167_));
 sky130_fd_sc_hd__o21ai_0 _25924_ (.A1(_10873_),
    .A2(_07166_),
    .B1(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__o211ai_1 _25925_ (.A1(_10898_),
    .A2(_07160_),
    .B1(_07163_),
    .C1(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__o221ai_2 _25926_ (.A1(_07137_),
    .A2(_07148_),
    .B1(_07153_),
    .B2(_07158_),
    .C1(_07169_),
    .Y(\if_stage_i.compressed_decoder_i.illegal_instr_o ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_59 ();
 sky130_fd_sc_hd__o21ai_2 _25929_ (.A1(_10776_),
    .A2(_07140_),
    .B1(net3733),
    .Y(_07172_));
 sky130_fd_sc_hd__nand2_1 _25930_ (.A(_10767_),
    .B(_07172_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[0] ));
 sky130_fd_sc_hd__nor4_2 _25931_ (.A(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .B(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .C(_10892_),
    .D(_07145_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand3_1 _25932_ (.A(_10767_),
    .B(_07173_),
    .C(_07141_),
    .Y(_07174_));
 sky130_fd_sc_hd__o21ai_0 _25933_ (.A1(_10767_),
    .A2(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .B1(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_58 ();
 sky130_fd_sc_hd__o21ai_0 _25935_ (.A1(_10769_),
    .A2(_10878_),
    .B1(_10775_),
    .Y(_07177_));
 sky130_fd_sc_hd__a21oi_1 _25936_ (.A1(_10769_),
    .A2(_07140_),
    .B1(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__nor2_1 _25937_ (.A(_10776_),
    .B(_10873_),
    .Y(_07179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__a21oi_1 _25939_ (.A1(_10769_),
    .A2(_07179_),
    .B1(_10858_),
    .Y(_07181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__o22ai_1 _25941_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .A2(_07178_),
    .B1(_07181_),
    .B2(_10866_),
    .Y(_07183_));
 sky130_fd_sc_hd__a21oi_1 _25942_ (.A1(_10776_),
    .A2(_07175_),
    .B1(_07183_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[10] ));
 sky130_fd_sc_hd__nand2_1 _25943_ (.A(_10776_),
    .B(_07174_),
    .Y(_07184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__nand2_4 _25945_ (.A(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .B(_10862_),
    .Y(_07186_));
 sky130_fd_sc_hd__nor2_4 _25946_ (.A(_10896_),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__nand2_2 _25947_ (.A(_07141_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__a31oi_1 _25948_ (.A1(_10872_),
    .A2(_07157_),
    .A3(_07188_),
    .B1(_10767_),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_1 _25949_ (.A(_10769_),
    .B(_07159_),
    .Y(_07190_));
 sky130_fd_sc_hd__o21ai_0 _25950_ (.A1(_07189_),
    .A2(_07190_),
    .B1(_10775_),
    .Y(_07191_));
 sky130_fd_sc_hd__a21boi_0 _25951_ (.A1(_07184_),
    .A2(_07191_),
    .B1_N(_10862_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[11] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__nand2_4 _25953_ (.A(_10767_),
    .B(_10776_),
    .Y(_07193_));
 sky130_fd_sc_hd__nor2_4 _25954_ (.A(_10767_),
    .B(_10775_),
    .Y(_07194_));
 sky130_fd_sc_hd__a31oi_2 _25955_ (.A1(_07157_),
    .A2(_07150_),
    .A3(_07151_),
    .B1(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__o21ai_2 _25956_ (.A1(_10866_),
    .A2(_07193_),
    .B1(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__clkinv_1 _25957_ (.A(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__nor2_4 _25958_ (.A(_10873_),
    .B(_07157_),
    .Y(_07198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__nand3_2 _25960_ (.A(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .B(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .C(_10896_),
    .Y(_07200_));
 sky130_fd_sc_hd__nand2_1 _25961_ (.A(_10896_),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__o21ai_0 _25962_ (.A1(_07186_),
    .A2(_07201_),
    .B1(_07141_),
    .Y(_07202_));
 sky130_fd_sc_hd__nor2_4 _25963_ (.A(_10872_),
    .B(_10878_),
    .Y(_07203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__nand2_2 _25965_ (.A(_10850_),
    .B(_07154_),
    .Y(_07205_));
 sky130_fd_sc_hd__and2_4 _25966_ (.A(_07143_),
    .B(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__nand2_4 _25967_ (.A(_10867_),
    .B(_10872_),
    .Y(_07207_));
 sky130_fd_sc_hd__nor2_4 _25968_ (.A(_10896_),
    .B(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__a221oi_1 _25969_ (.A1(_10867_),
    .A2(_07203_),
    .B1(_07206_),
    .B2(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .C1(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__a21oi_1 _25970_ (.A1(_07202_),
    .A2(_07209_),
    .B1(_07137_),
    .Y(_07210_));
 sky130_fd_sc_hd__a21oi_1 _25971_ (.A1(_07163_),
    .A2(_07198_),
    .B1(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_2 _25972_ (.A1(_10896_),
    .A2(_07197_),
    .B1(_07211_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[12] ));
 sky130_fd_sc_hd__nor2_1 _25973_ (.A(_10838_),
    .B(_10898_),
    .Y(_07212_));
 sky130_fd_sc_hd__nor2_4 _25974_ (.A(_10873_),
    .B(_10878_),
    .Y(_07213_));
 sky130_fd_sc_hd__o2111ai_1 _25975_ (.A1(_10858_),
    .A2(_07212_),
    .B1(_07213_),
    .C1(net3733),
    .D1(_10862_),
    .Y(_07214_));
 sky130_fd_sc_hd__o21ai_1 _25976_ (.A1(_10896_),
    .A2(_07207_),
    .B1(_10775_),
    .Y(_07215_));
 sky130_fd_sc_hd__a31oi_1 _25977_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .A2(_07143_),
    .A3(_07205_),
    .B1(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__nand2_1 _25978_ (.A(_07214_),
    .B(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__o21ai_2 _25979_ (.A1(_10775_),
    .A2(_10867_),
    .B1(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__nand2_2 _25980_ (.A(_10866_),
    .B(_10872_),
    .Y(_07219_));
 sky130_fd_sc_hd__a21oi_1 _25981_ (.A1(_10769_),
    .A2(_10879_),
    .B1(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__a21oi_2 _25982_ (.A1(_10769_),
    .A2(_07218_),
    .B1(_07220_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[13] ));
 sky130_fd_sc_hd__nand2_8 _25983_ (.A(net3733),
    .B(_07213_),
    .Y(_07221_));
 sky130_fd_sc_hd__a21oi_1 _25984_ (.A1(_10896_),
    .A2(_07145_),
    .B1(_07186_),
    .Y(_07222_));
 sky130_fd_sc_hd__nor2_1 _25985_ (.A(_07221_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__a211oi_1 _25986_ (.A1(_10892_),
    .A2(_07206_),
    .B1(_07215_),
    .C1(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__a21oi_1 _25987_ (.A1(_10775_),
    .A2(_07157_),
    .B1(_10873_),
    .Y(_07225_));
 sky130_fd_sc_hd__nand3_1 _25988_ (.A(_10767_),
    .B(_10867_),
    .C(_10873_),
    .Y(_07226_));
 sky130_fd_sc_hd__o31ai_1 _25989_ (.A1(_10767_),
    .A2(_07224_),
    .A3(_07225_),
    .B1(_07226_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[14] ));
 sky130_fd_sc_hd__nor2_2 _25990_ (.A(_07156_),
    .B(_07221_),
    .Y(_07227_));
 sky130_fd_sc_hd__and2_4 _25991_ (.A(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .B(_10862_),
    .X(_07228_));
 sky130_fd_sc_hd__nand2_4 _25992_ (.A(_10898_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__o21ai_0 _25993_ (.A1(_10846_),
    .A2(_07200_),
    .B1(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__nand2_2 _25994_ (.A(_07228_),
    .B(_07201_),
    .Y(_07231_));
 sky130_fd_sc_hd__nand2_4 _25995_ (.A(_07141_),
    .B(_07231_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_1 _25996_ (.A(_10873_),
    .B(_10879_),
    .Y(_07233_));
 sky130_fd_sc_hd__a21oi_1 _25997_ (.A1(_07160_),
    .A2(_07233_),
    .B1(_10846_),
    .Y(_07234_));
 sky130_fd_sc_hd__a211oi_1 _25998_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .A2(_07206_),
    .B1(_07234_),
    .C1(_07208_),
    .Y(_07235_));
 sky130_fd_sc_hd__o21ai_0 _25999_ (.A1(_10846_),
    .A2(_07232_),
    .B1(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__a21oi_1 _26000_ (.A1(_07227_),
    .A2(_07230_),
    .B1(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__nor2_1 _26001_ (.A(_07137_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__a21oi_1 _26002_ (.A1(_10867_),
    .A2(_10879_),
    .B1(_07198_),
    .Y(_07239_));
 sky130_fd_sc_hd__nand2_2 _26003_ (.A(_10896_),
    .B(_07146_),
    .Y(_07240_));
 sky130_fd_sc_hd__nand2_2 _26004_ (.A(_07141_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a21oi_1 _26005_ (.A1(_07239_),
    .A2(_07241_),
    .B1(_07193_),
    .Y(_07242_));
 sky130_fd_sc_hd__nor2b_1 _26006_ (.A(_07238_),
    .B_N(_07239_),
    .Y(_07243_));
 sky130_fd_sc_hd__o21ai_0 _26007_ (.A1(_07198_),
    .A2(_07243_),
    .B1(_10846_),
    .Y(_07244_));
 sky130_fd_sc_hd__o21ai_0 _26008_ (.A1(_07238_),
    .A2(_07242_),
    .B1(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__nor2_1 _26009_ (.A(_10846_),
    .B(_07150_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21oi_1 _26010_ (.A1(_10879_),
    .A2(_07150_),
    .B1(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__nand2_8 _26011_ (.A(_10767_),
    .B(_10775_),
    .Y(_07248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__o21ai_0 _26013_ (.A1(_10775_),
    .A2(_10878_),
    .B1(_07245_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_1 _26014_ (.A(_10769_),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__o221ai_1 _26015_ (.A1(_10775_),
    .A2(_07245_),
    .B1(_07247_),
    .B2(_07248_),
    .C1(_07251_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[15] ));
 sky130_fd_sc_hd__mux2_8 _26016_ (.A0(_10765_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ),
    .S(net3948),
    .X(_07252_));
 sky130_fd_sc_hd__o21ai_0 _26017_ (.A1(_10866_),
    .A2(_07252_),
    .B1(_07163_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21oi_1 _26018_ (.A1(_10850_),
    .A2(_07240_),
    .B1(_07221_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_1 _26019_ (.A(_10850_),
    .B(_10873_),
    .Y(_07255_));
 sky130_fd_sc_hd__a21oi_1 _26020_ (.A1(_10867_),
    .A2(_07154_),
    .B1(_10879_),
    .Y(_07256_));
 sky130_fd_sc_hd__nor3_1 _26021_ (.A(_10838_),
    .B(_10872_),
    .C(_10879_),
    .Y(_07257_));
 sky130_fd_sc_hd__a21oi_1 _26022_ (.A1(_10872_),
    .A2(_10898_),
    .B1(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__o22ai_1 _26023_ (.A1(_07255_),
    .A2(_07256_),
    .B1(_07258_),
    .B2(_10866_),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_1 _26024_ (.A(_10850_),
    .B(_07229_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _26025_ (.A(_07187_),
    .B(_07252_),
    .Y(_07261_));
 sky130_fd_sc_hd__a31oi_1 _26026_ (.A1(_10879_),
    .A2(_07260_),
    .A3(_07261_),
    .B1(_07219_),
    .Y(_07262_));
 sky130_fd_sc_hd__nor2_4 _26027_ (.A(_10767_),
    .B(_10776_),
    .Y(_07263_));
 sky130_fd_sc_hd__o21ai_0 _26028_ (.A1(_07259_),
    .A2(_07262_),
    .B1(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__o21ai_0 _26029_ (.A1(_07253_),
    .A2(_07254_),
    .B1(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__o21ai_0 _26030_ (.A1(_10850_),
    .A2(_07160_),
    .B1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_1 _26031_ (.A(_10776_),
    .B(_07252_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_1 _26032_ (.A(_10769_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand2_1 _26033_ (.A(_07193_),
    .B(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__nor2_4 _26034_ (.A(_10867_),
    .B(_10872_),
    .Y(_07270_));
 sky130_fd_sc_hd__nand2_8 _26035_ (.A(_10866_),
    .B(_07140_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_1 _26036_ (.A(_07160_),
    .B(_07151_),
    .Y(_07272_));
 sky130_fd_sc_hd__a221oi_1 _26037_ (.A1(_10850_),
    .A2(_07270_),
    .B1(_07252_),
    .B2(_07271_),
    .C1(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__a21oi_1 _26038_ (.A1(_07266_),
    .A2(_07269_),
    .B1(_07273_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[16] ));
 sky130_fd_sc_hd__nand2_2 _26039_ (.A(net3948),
    .B(_10900_),
    .Y(_07274_));
 sky130_fd_sc_hd__o21ai_4 _26040_ (.A1(net3948),
    .A2(_10773_),
    .B1(_07274_),
    .Y(_07275_));
 sky130_fd_sc_hd__o221ai_1 _26041_ (.A1(_10854_),
    .A2(_07241_),
    .B1(_07275_),
    .B2(_10866_),
    .C1(_07160_),
    .Y(_07276_));
 sky130_fd_sc_hd__a21oi_1 _26042_ (.A1(_07141_),
    .A2(_07229_),
    .B1(_07203_),
    .Y(_07277_));
 sky130_fd_sc_hd__and3_4 _26043_ (.A(_10898_),
    .B(_07143_),
    .C(_07205_),
    .X(_07278_));
 sky130_fd_sc_hd__nor3_2 _26044_ (.A(_07198_),
    .B(_07208_),
    .C(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__o221ai_1 _26045_ (.A1(_07188_),
    .A2(_07275_),
    .B1(_07277_),
    .B2(_10854_),
    .C1(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__a22o_1 _26046_ (.A1(_07163_),
    .A2(_07276_),
    .B1(_07280_),
    .B2(_07263_),
    .X(_07281_));
 sky130_fd_sc_hd__a31oi_1 _26047_ (.A1(_10866_),
    .A2(_10873_),
    .A3(_07151_),
    .B1(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__nand2_1 _26048_ (.A(_07160_),
    .B(_07281_),
    .Y(_07283_));
 sky130_fd_sc_hd__o221ai_1 _26049_ (.A1(_07195_),
    .A2(_07275_),
    .B1(_07282_),
    .B2(_10854_),
    .C1(_07283_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[17] ));
 sky130_fd_sc_hd__nand2_1 _26050_ (.A(net3948),
    .B(_10901_),
    .Y(_07284_));
 sky130_fd_sc_hd__o21ai_4 _26051_ (.A1(net3948),
    .A2(_10886_),
    .B1(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__o221ai_1 _26052_ (.A1(_10858_),
    .A2(_07241_),
    .B1(_07285_),
    .B2(_10866_),
    .C1(_07160_),
    .Y(_07286_));
 sky130_fd_sc_hd__nand2_4 _26053_ (.A(net3733),
    .B(_10879_),
    .Y(_07287_));
 sky130_fd_sc_hd__a21oi_1 _26054_ (.A1(_07187_),
    .A2(_07285_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nor2_1 _26055_ (.A(_07203_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__a21oi_1 _26056_ (.A1(_07279_),
    .A2(_07289_),
    .B1(_07137_),
    .Y(_07290_));
 sky130_fd_sc_hd__a21oi_1 _26057_ (.A1(_07163_),
    .A2(_07286_),
    .B1(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__a21oi_1 _26058_ (.A1(_10858_),
    .A2(_07198_),
    .B1(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__o21ai_0 _26059_ (.A1(_07159_),
    .A2(_07285_),
    .B1(_07150_),
    .Y(_07293_));
 sky130_fd_sc_hd__a22oi_1 _26060_ (.A1(_10776_),
    .A2(_07292_),
    .B1(_07293_),
    .B2(_07151_),
    .Y(_07294_));
 sky130_fd_sc_hd__nor2_1 _26061_ (.A(_10775_),
    .B(_07285_),
    .Y(_07295_));
 sky130_fd_sc_hd__o21ai_0 _26062_ (.A1(_07292_),
    .A2(_07295_),
    .B1(_10769_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_1 _26063_ (.A(_07294_),
    .B(_07296_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[18] ));
 sky130_fd_sc_hd__mux2i_2 _26064_ (.A0(_10882_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ),
    .S(net3948),
    .Y(_07297_));
 sky130_fd_sc_hd__a21oi_1 _26065_ (.A1(_10862_),
    .A2(_07240_),
    .B1(_10878_),
    .Y(_07298_));
 sky130_fd_sc_hd__o22ai_1 _26066_ (.A1(_10866_),
    .A2(_07297_),
    .B1(_07298_),
    .B2(_07219_),
    .Y(_07299_));
 sky130_fd_sc_hd__o21ai_0 _26067_ (.A1(_07188_),
    .A2(_07297_),
    .B1(_07279_),
    .Y(_07300_));
 sky130_fd_sc_hd__a22oi_1 _26068_ (.A1(_07163_),
    .A2(_07299_),
    .B1(_07300_),
    .B2(_07263_),
    .Y(_07301_));
 sky130_fd_sc_hd__nor2_1 _26069_ (.A(_10862_),
    .B(_07160_),
    .Y(_07302_));
 sky130_fd_sc_hd__o22ai_1 _26070_ (.A1(_07195_),
    .A2(_07297_),
    .B1(_07301_),
    .B2(_07302_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[19] ));
 sky130_fd_sc_hd__nor2_4 _26071_ (.A(_07221_),
    .B(_07229_),
    .Y(_07303_));
 sky130_fd_sc_hd__nor2_4 _26072_ (.A(_10867_),
    .B(_07213_),
    .Y(_07304_));
 sky130_fd_sc_hd__a21oi_1 _26073_ (.A1(_10767_),
    .A2(_07304_),
    .B1(_10776_),
    .Y(_07305_));
 sky130_fd_sc_hd__o21ai_2 _26074_ (.A1(_10767_),
    .A2(_07303_),
    .B1(_07305_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[1] ));
 sky130_fd_sc_hd__nand2_2 _26075_ (.A(_10898_),
    .B(_07155_),
    .Y(_07306_));
 sky130_fd_sc_hd__o21ai_0 _26076_ (.A1(_07146_),
    .A2(_07306_),
    .B1(_10888_),
    .Y(_07307_));
 sky130_fd_sc_hd__o21ai_0 _26077_ (.A1(_10878_),
    .A2(_10888_),
    .B1(_10873_),
    .Y(_07308_));
 sky130_fd_sc_hd__mux2i_4 _26078_ (.A0(_10890_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ),
    .S(net3948),
    .Y(_07309_));
 sky130_fd_sc_hd__nor2_1 _26079_ (.A(_10866_),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__a31oi_1 _26080_ (.A1(_10866_),
    .A2(_07307_),
    .A3(_07308_),
    .B1(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__o21ai_0 _26081_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .A2(_07160_),
    .B1(_07163_),
    .Y(_07312_));
 sky130_fd_sc_hd__nor2_4 _26082_ (.A(_07198_),
    .B(_07137_),
    .Y(_07313_));
 sky130_fd_sc_hd__o22ai_1 _26083_ (.A1(_10888_),
    .A2(_07200_),
    .B1(_07309_),
    .B2(_07229_),
    .Y(_07314_));
 sky130_fd_sc_hd__a211oi_1 _26084_ (.A1(_07227_),
    .A2(_07314_),
    .B1(_07278_),
    .C1(_07208_),
    .Y(_07315_));
 sky130_fd_sc_hd__o21ai_0 _26085_ (.A1(_10888_),
    .A2(_07232_),
    .B1(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nor2_1 _26086_ (.A(_10775_),
    .B(_07309_),
    .Y(_07317_));
 sky130_fd_sc_hd__a31oi_1 _26087_ (.A1(_10775_),
    .A2(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .A3(_07159_),
    .B1(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__o22ai_1 _26088_ (.A1(_10888_),
    .A2(_07150_),
    .B1(_07309_),
    .B2(_10873_),
    .Y(_07319_));
 sky130_fd_sc_hd__a21oi_1 _26089_ (.A1(_10879_),
    .A2(_07319_),
    .B1(_07310_),
    .Y(_07320_));
 sky130_fd_sc_hd__o22ai_1 _26090_ (.A1(_10767_),
    .A2(_07318_),
    .B1(_07320_),
    .B2(_07248_),
    .Y(_07321_));
 sky130_fd_sc_hd__a21oi_1 _26091_ (.A1(_07313_),
    .A2(_07316_),
    .B1(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__o21ai_0 _26092_ (.A1(_07311_),
    .A2(_07312_),
    .B1(_07322_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[20] ));
 sky130_fd_sc_hd__mux2i_2 _26093_ (.A0(_10840_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .S(net3948),
    .Y(_07323_));
 sky130_fd_sc_hd__nor2_4 _26094_ (.A(_10872_),
    .B(_10879_),
    .Y(_07324_));
 sky130_fd_sc_hd__nor2_1 _26095_ (.A(_07140_),
    .B(_07200_),
    .Y(_07325_));
 sky130_fd_sc_hd__o21ai_2 _26096_ (.A1(_07324_),
    .A2(_07325_),
    .B1(_10866_),
    .Y(_07326_));
 sky130_fd_sc_hd__nand2_2 _26097_ (.A(_10898_),
    .B(_07206_),
    .Y(_07327_));
 sky130_fd_sc_hd__o221ai_1 _26098_ (.A1(_07188_),
    .A2(_07323_),
    .B1(_07326_),
    .B2(_10884_),
    .C1(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nand2_1 _26099_ (.A(_07313_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__nor2_2 _26100_ (.A(_10769_),
    .B(_10867_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand3_1 _26101_ (.A(_10767_),
    .B(_10879_),
    .C(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .Y(_07331_));
 sky130_fd_sc_hd__o22ai_1 _26102_ (.A1(_07323_),
    .A2(_07330_),
    .B1(_07331_),
    .B2(_07150_),
    .Y(_07332_));
 sky130_fd_sc_hd__a22oi_1 _26103_ (.A1(_10866_),
    .A2(_07163_),
    .B1(_07263_),
    .B2(_07287_),
    .Y(_07333_));
 sky130_fd_sc_hd__o22ai_1 _26104_ (.A1(_07137_),
    .A2(_07232_),
    .B1(_07333_),
    .B2(_10873_),
    .Y(_07334_));
 sky130_fd_sc_hd__nor2_1 _26105_ (.A(_10873_),
    .B(_07323_),
    .Y(_07335_));
 sky130_fd_sc_hd__a21oi_1 _26106_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .A2(_07270_),
    .B1(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__o22ai_1 _26107_ (.A1(_10866_),
    .A2(_07323_),
    .B1(_07336_),
    .B2(_10878_),
    .Y(_07337_));
 sky130_fd_sc_hd__a222oi_1 _26108_ (.A1(_10776_),
    .A2(_07332_),
    .B1(_07334_),
    .B2(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .C1(_07151_),
    .C2(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_2 _26109_ (.A(_07329_),
    .B(_07338_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[21] ));
 sky130_fd_sc_hd__nand2_1 _26110_ (.A(_10892_),
    .B(_07203_),
    .Y(_07339_));
 sky130_fd_sc_hd__o21ai_0 _26111_ (.A1(_10838_),
    .A2(_10879_),
    .B1(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nor2_1 _26112_ (.A(net3948),
    .B(_10833_),
    .Y(_07341_));
 sky130_fd_sc_hd__a21oi_2 _26113_ (.A1(net3948),
    .A2(_10903_),
    .B1(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__a221oi_1 _26114_ (.A1(_10866_),
    .A2(_07340_),
    .B1(_07342_),
    .B2(_07271_),
    .C1(_07248_),
    .Y(_07343_));
 sky130_fd_sc_hd__nand2_1 _26115_ (.A(_07232_),
    .B(_07326_),
    .Y(_07344_));
 sky130_fd_sc_hd__a221o_1 _26116_ (.A1(_07303_),
    .A2(_07342_),
    .B1(_07344_),
    .B2(_10892_),
    .C1(_07278_),
    .X(_07345_));
 sky130_fd_sc_hd__nand3_1 _26117_ (.A(_10769_),
    .B(_07179_),
    .C(_07287_),
    .Y(_07346_));
 sky130_fd_sc_hd__o41ai_1 _26118_ (.A1(_10769_),
    .A2(_10775_),
    .A3(_10867_),
    .A4(_07203_),
    .B1(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a31oi_1 _26119_ (.A1(_10879_),
    .A2(_10892_),
    .A3(_07270_),
    .B1(_10775_),
    .Y(_07348_));
 sky130_fd_sc_hd__a21oi_1 _26120_ (.A1(_10767_),
    .A2(_10867_),
    .B1(_07194_),
    .Y(_07349_));
 sky130_fd_sc_hd__inv_1 _26121_ (.A(_07342_),
    .Y(_07350_));
 sky130_fd_sc_hd__o22ai_1 _26122_ (.A1(_10769_),
    .A2(_07348_),
    .B1(_07349_),
    .B2(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__a221oi_1 _26123_ (.A1(_07313_),
    .A2(_07345_),
    .B1(_07347_),
    .B2(_10892_),
    .C1(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__nor2_2 _26124_ (.A(_07343_),
    .B(_07352_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[22] ));
 sky130_fd_sc_hd__nor2_1 _26125_ (.A(net3948),
    .B(_10844_),
    .Y(_07353_));
 sky130_fd_sc_hd__a21oi_2 _26126_ (.A1(net3948),
    .A2(_10904_),
    .B1(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__nor2_1 _26127_ (.A(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .B(_10873_),
    .Y(_07355_));
 sky130_fd_sc_hd__a21oi_1 _26128_ (.A1(_10858_),
    .A2(_10873_),
    .B1(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__o22ai_2 _26129_ (.A1(_07304_),
    .A2(_07354_),
    .B1(_07356_),
    .B2(_07157_),
    .Y(_07357_));
 sky130_fd_sc_hd__nor2_2 _26130_ (.A(_10842_),
    .B(_07150_),
    .Y(_07358_));
 sky130_fd_sc_hd__o21ai_0 _26131_ (.A1(_10896_),
    .A2(_07354_),
    .B1(_07228_),
    .Y(_07359_));
 sky130_fd_sc_hd__o21ai_0 _26132_ (.A1(_10842_),
    .A2(_07228_),
    .B1(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__a221oi_1 _26133_ (.A1(_10878_),
    .A2(_07358_),
    .B1(_07360_),
    .B2(_07141_),
    .C1(_07278_),
    .Y(_07361_));
 sky130_fd_sc_hd__a21oi_1 _26134_ (.A1(_10879_),
    .A2(_07358_),
    .B1(_10775_),
    .Y(_07362_));
 sky130_fd_sc_hd__nor2_1 _26135_ (.A(_10769_),
    .B(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__a21oi_1 _26136_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .A2(_07347_),
    .B1(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__nand2b_1 _26137_ (.A_N(_07349_),
    .B(_07354_),
    .Y(_07365_));
 sky130_fd_sc_hd__o311a_4 _26138_ (.A1(_07198_),
    .A2(_07137_),
    .A3(_07361_),
    .B1(_07364_),
    .C1(_07365_),
    .X(_07366_));
 sky130_fd_sc_hd__a21oi_4 _26139_ (.A1(_07151_),
    .A2(_07357_),
    .B1(_07366_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[23] ));
 sky130_fd_sc_hd__mux2_8 _26140_ (.A0(_10848_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .S(net3948),
    .X(_07367_));
 sky130_fd_sc_hd__nor2_1 _26141_ (.A(_10873_),
    .B(_10879_),
    .Y(_07368_));
 sky130_fd_sc_hd__and3_4 _26142_ (.A(_10850_),
    .B(_07154_),
    .C(_07143_),
    .X(_07369_));
 sky130_fd_sc_hd__a21oi_2 _26143_ (.A1(_07141_),
    .A2(_07186_),
    .B1(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__nor2_4 _26144_ (.A(_10866_),
    .B(_10873_),
    .Y(_07371_));
 sky130_fd_sc_hd__a21oi_1 _26145_ (.A1(_10838_),
    .A2(_10873_),
    .B1(_07157_),
    .Y(_07372_));
 sky130_fd_sc_hd__a221oi_1 _26146_ (.A1(_10862_),
    .A2(_07371_),
    .B1(_07367_),
    .B2(_07303_),
    .C1(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__o211ai_1 _26147_ (.A1(_10838_),
    .A2(_07370_),
    .B1(_07373_),
    .C1(_07327_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2_1 _26148_ (.A(_07263_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__o211ai_1 _26149_ (.A1(_07368_),
    .A2(_07375_),
    .B1(_10838_),
    .C1(_10866_),
    .Y(_07376_));
 sky130_fd_sc_hd__o21ai_0 _26150_ (.A1(_10866_),
    .A2(_07367_),
    .B1(_07163_),
    .Y(_07377_));
 sky130_fd_sc_hd__nand2_1 _26151_ (.A(_07375_),
    .B(_07377_),
    .Y(_07378_));
 sky130_fd_sc_hd__a221oi_1 _26152_ (.A1(_07194_),
    .A2(_07367_),
    .B1(_07376_),
    .B2(_07378_),
    .C1(_07151_),
    .Y(_07379_));
 sky130_fd_sc_hd__a221oi_1 _26153_ (.A1(_10862_),
    .A2(_07159_),
    .B1(_07271_),
    .B2(_07367_),
    .C1(_07248_),
    .Y(_07380_));
 sky130_fd_sc_hd__nor2_1 _26154_ (.A(_07379_),
    .B(_07380_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[24] ));
 sky130_fd_sc_hd__nor2_1 _26155_ (.A(net3948),
    .B(_10852_),
    .Y(_07381_));
 sky130_fd_sc_hd__a21oi_2 _26156_ (.A1(net3948),
    .A2(_10905_),
    .B1(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__nor2_1 _26157_ (.A(_10896_),
    .B(_07271_),
    .Y(_07383_));
 sky130_fd_sc_hd__a21oi_1 _26158_ (.A1(_07271_),
    .A2(_07382_),
    .B1(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__nor2_2 _26159_ (.A(_10872_),
    .B(_10896_),
    .Y(_07385_));
 sky130_fd_sc_hd__mux2i_1 _26160_ (.A0(_07382_),
    .A1(_07385_),
    .S(_07330_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21oi_1 _26161_ (.A1(_10873_),
    .A2(_07205_),
    .B1(_10866_),
    .Y(_07387_));
 sky130_fd_sc_hd__a211oi_2 _26162_ (.A1(_10873_),
    .A2(_10896_),
    .B1(_07387_),
    .C1(_10879_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand3_4 _26163_ (.A(_10862_),
    .B(_10898_),
    .C(_07141_),
    .Y(_07389_));
 sky130_fd_sc_hd__nor2_1 _26164_ (.A(_10858_),
    .B(_07382_),
    .Y(_07390_));
 sky130_fd_sc_hd__nor2_1 _26165_ (.A(_07389_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nor3_1 _26166_ (.A(_07371_),
    .B(_07203_),
    .C(_07369_),
    .Y(_07392_));
 sky130_fd_sc_hd__nor2_1 _26167_ (.A(_10888_),
    .B(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__a21oi_4 _26168_ (.A1(_10896_),
    .A2(_07198_),
    .B1(_07137_),
    .Y(_07394_));
 sky130_fd_sc_hd__o31ai_1 _26169_ (.A1(_07388_),
    .A2(_07391_),
    .A3(_07393_),
    .B1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__o221ai_2 _26170_ (.A1(_07248_),
    .A2(_07384_),
    .B1(_07386_),
    .B2(_10775_),
    .C1(_07395_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[25] ));
 sky130_fd_sc_hd__nor2_1 _26171_ (.A(net3948),
    .B(_10856_),
    .Y(_07396_));
 sky130_fd_sc_hd__a21oi_2 _26172_ (.A1(net3948),
    .A2(_10906_),
    .B1(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__nor2_1 _26173_ (.A(_10858_),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__o21ai_0 _26174_ (.A1(_07203_),
    .A2(_07369_),
    .B1(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .Y(_07399_));
 sky130_fd_sc_hd__o221ai_1 _26175_ (.A1(_10846_),
    .A2(_07207_),
    .B1(_07389_),
    .B2(_07398_),
    .C1(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__o21ai_0 _26176_ (.A1(_07388_),
    .A2(_07400_),
    .B1(_07394_),
    .Y(_07401_));
 sky130_fd_sc_hd__nand2_1 _26177_ (.A(\if_stage_i.compressed_decoder_i.instr_i[7] ),
    .B(_10879_),
    .Y(_07402_));
 sky130_fd_sc_hd__o21ai_0 _26178_ (.A1(_10879_),
    .A2(_10888_),
    .B1(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__nor2_1 _26179_ (.A(_10775_),
    .B(_07330_),
    .Y(_07404_));
 sky130_fd_sc_hd__a32oi_1 _26180_ (.A1(_07163_),
    .A2(_07270_),
    .A3(_07403_),
    .B1(_07404_),
    .B2(_07397_),
    .Y(_07405_));
 sky130_fd_sc_hd__nor2_1 _26181_ (.A(_10846_),
    .B(_07160_),
    .Y(_07406_));
 sky130_fd_sc_hd__a2111oi_0 _26182_ (.A1(_07271_),
    .A2(_07397_),
    .B1(_07406_),
    .C1(_07358_),
    .D1(_07248_),
    .Y(_07407_));
 sky130_fd_sc_hd__a31oi_2 _26183_ (.A1(_07248_),
    .A2(_07401_),
    .A3(_07405_),
    .B1(_07407_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[26] ));
 sky130_fd_sc_hd__nand2_1 _26184_ (.A(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .B(_07143_),
    .Y(_07408_));
 sky130_fd_sc_hd__nor2_4 _26185_ (.A(_07371_),
    .B(_07203_),
    .Y(_07409_));
 sky130_fd_sc_hd__o22ai_1 _26186_ (.A1(_07205_),
    .A2(_07408_),
    .B1(_07409_),
    .B2(_10838_),
    .Y(_07410_));
 sky130_fd_sc_hd__nand2_1 _26187_ (.A(net3948),
    .B(_10907_),
    .Y(_07411_));
 sky130_fd_sc_hd__o21ai_2 _26188_ (.A1(net3948),
    .A2(_10860_),
    .B1(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__a21oi_1 _26189_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .A2(_07412_),
    .B1(_07389_),
    .Y(_07413_));
 sky130_fd_sc_hd__o31ai_1 _26190_ (.A1(_07388_),
    .A2(_07410_),
    .A3(_07413_),
    .B1(_07394_),
    .Y(_07414_));
 sky130_fd_sc_hd__nor2_1 _26191_ (.A(_10879_),
    .B(_10884_),
    .Y(_07415_));
 sky130_fd_sc_hd__a21oi_1 _26192_ (.A1(_10850_),
    .A2(_10879_),
    .B1(_07415_),
    .Y(_07416_));
 sky130_fd_sc_hd__o21ai_0 _26193_ (.A1(_10769_),
    .A2(_10867_),
    .B1(_10776_),
    .Y(_07417_));
 sky130_fd_sc_hd__o32a_1 _26194_ (.A1(_07193_),
    .A2(_07150_),
    .A3(_07416_),
    .B1(_07412_),
    .B2(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__nor2_1 _26195_ (.A(_07304_),
    .B(_07412_),
    .Y(_07419_));
 sky130_fd_sc_hd__a211oi_1 _26196_ (.A1(_10850_),
    .A2(_07198_),
    .B1(_07248_),
    .C1(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__a31oi_2 _26197_ (.A1(_07248_),
    .A2(_07414_),
    .A3(_07418_),
    .B1(_07420_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[27] ));
 sky130_fd_sc_hd__mux2_8 _26198_ (.A0(_10894_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ),
    .S(net3948),
    .X(_07421_));
 sky130_fd_sc_hd__a221oi_1 _26199_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .A2(_07198_),
    .B1(_07271_),
    .B2(_07421_),
    .C1(_07248_),
    .Y(_07422_));
 sky130_fd_sc_hd__nor2_1 _26200_ (.A(_10858_),
    .B(_07421_),
    .Y(_07423_));
 sky130_fd_sc_hd__nand2_1 _26201_ (.A(_10892_),
    .B(_07369_),
    .Y(_07424_));
 sky130_fd_sc_hd__nor2_1 _26202_ (.A(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .B(_10873_),
    .Y(_07425_));
 sky130_fd_sc_hd__o21ai_0 _26203_ (.A1(_07324_),
    .A2(_07425_),
    .B1(_10867_),
    .Y(_07426_));
 sky130_fd_sc_hd__a21oi_1 _26204_ (.A1(_10873_),
    .A2(_10896_),
    .B1(_07141_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21oi_1 _26205_ (.A1(_07426_),
    .A2(_07427_),
    .B1(_07278_),
    .Y(_07428_));
 sky130_fd_sc_hd__o211ai_1 _26206_ (.A1(_07389_),
    .A2(_07423_),
    .B1(_07424_),
    .C1(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__a221oi_2 _26207_ (.A1(_07404_),
    .A2(_07421_),
    .B1(_07429_),
    .B2(_07394_),
    .C1(_07151_),
    .Y(_07430_));
 sky130_fd_sc_hd__nor2_4 _26208_ (.A(_07422_),
    .B(_07430_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[28] ));
 sky130_fd_sc_hd__a21oi_1 _26209_ (.A1(_10858_),
    .A2(_10867_),
    .B1(_10873_),
    .Y(_07431_));
 sky130_fd_sc_hd__mux2i_2 _26210_ (.A0(_10864_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ),
    .S(net3948),
    .Y(_07432_));
 sky130_fd_sc_hd__a21oi_1 _26211_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .A2(_07432_),
    .B1(_07389_),
    .Y(_07433_));
 sky130_fd_sc_hd__a211o_1 _26212_ (.A1(_07287_),
    .A2(_07431_),
    .B1(_07433_),
    .C1(_07385_),
    .X(_07434_));
 sky130_fd_sc_hd__o22ai_1 _26213_ (.A1(_10858_),
    .A2(_07160_),
    .B1(_07304_),
    .B2(_07432_),
    .Y(_07435_));
 sky130_fd_sc_hd__nor2_1 _26214_ (.A(_07417_),
    .B(_07432_),
    .Y(_07436_));
 sky130_fd_sc_hd__a221o_1 _26215_ (.A1(_07394_),
    .A2(_07434_),
    .B1(_07435_),
    .B2(_07151_),
    .C1(_07436_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[29] ));
 sky130_fd_sc_hd__o22ai_2 _26216_ (.A1(_10769_),
    .A2(_07172_),
    .B1(_07303_),
    .B2(_07137_),
    .Y(_07437_));
 sky130_fd_sc_hd__o21ai_1 _26217_ (.A1(_07371_),
    .A2(_07206_),
    .B1(_07263_),
    .Y(_07438_));
 sky130_fd_sc_hd__nand4_1 _26218_ (.A(_07173_),
    .B(_07163_),
    .C(_07141_),
    .D(_07306_),
    .Y(_07439_));
 sky130_fd_sc_hd__o211ai_1 _26219_ (.A1(_10888_),
    .A2(_07437_),
    .B1(_07438_),
    .C1(_07439_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[2] ));
 sky130_fd_sc_hd__mux2i_1 _26220_ (.A0(_10870_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ),
    .S(net3948),
    .Y(_07440_));
 sky130_fd_sc_hd__o21ai_0 _26221_ (.A1(_10858_),
    .A2(_07440_),
    .B1(_07139_),
    .Y(_07441_));
 sky130_fd_sc_hd__nand3_1 _26222_ (.A(_10838_),
    .B(_10842_),
    .C(_10896_),
    .Y(_07442_));
 sky130_fd_sc_hd__a21oi_1 _26223_ (.A1(_10862_),
    .A2(_07442_),
    .B1(_10858_),
    .Y(_07443_));
 sky130_fd_sc_hd__a211oi_1 _26224_ (.A1(_10898_),
    .A2(_07441_),
    .B1(_07443_),
    .C1(_07287_),
    .Y(_07444_));
 sky130_fd_sc_hd__o21ai_0 _26225_ (.A1(_10850_),
    .A2(net3733),
    .B1(_10872_),
    .Y(_07445_));
 sky130_fd_sc_hd__nor2_1 _26226_ (.A(_07444_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__o21ai_0 _26227_ (.A1(_07385_),
    .A2(_07446_),
    .B1(_07394_),
    .Y(_07447_));
 sky130_fd_sc_hd__o21ai_0 _26228_ (.A1(_07197_),
    .A2(_07440_),
    .B1(_07447_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[30] ));
 sky130_fd_sc_hd__mux2_8 _26229_ (.A0(_10876_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .S(net3948),
    .X(_07448_));
 sky130_fd_sc_hd__o21ai_0 _26230_ (.A1(_10858_),
    .A2(_07448_),
    .B1(_10862_),
    .Y(_07449_));
 sky130_fd_sc_hd__nand2_1 _26231_ (.A(_07141_),
    .B(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__a32o_4 _26232_ (.A1(_10898_),
    .A2(_07263_),
    .A3(_07450_),
    .B1(_07448_),
    .B2(_07196_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[31] ));
 sky130_fd_sc_hd__o22ai_1 _26233_ (.A1(_07137_),
    .A2(_07207_),
    .B1(_07437_),
    .B2(_10884_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[3] ));
 sky130_fd_sc_hd__o21ai_0 _26234_ (.A1(_10892_),
    .A2(_07159_),
    .B1(_07150_),
    .Y(_07451_));
 sky130_fd_sc_hd__a21oi_1 _26235_ (.A1(_10879_),
    .A2(_07187_),
    .B1(_10776_),
    .Y(_07452_));
 sky130_fd_sc_hd__o22ai_1 _26236_ (.A1(_10776_),
    .A2(_07409_),
    .B1(_07452_),
    .B2(_10892_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21oi_1 _26237_ (.A1(_07173_),
    .A2(_07306_),
    .B1(_07221_),
    .Y(_07454_));
 sky130_fd_sc_hd__a2111oi_0 _26238_ (.A1(_10867_),
    .A2(_10892_),
    .B1(_07198_),
    .C1(_07454_),
    .D1(_10769_),
    .Y(_07455_));
 sky130_fd_sc_hd__a21oi_1 _26239_ (.A1(_10769_),
    .A2(_07453_),
    .B1(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__nor2_1 _26240_ (.A(_07151_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__a21oi_1 _26241_ (.A1(_07151_),
    .A2(_07451_),
    .B1(_07457_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[4] ));
 sky130_fd_sc_hd__o21ai_0 _26242_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .A2(_10896_),
    .B1(_07228_),
    .Y(_07458_));
 sky130_fd_sc_hd__o21ai_0 _26243_ (.A1(_10878_),
    .A2(_07458_),
    .B1(_07409_),
    .Y(_07459_));
 sky130_fd_sc_hd__o21ai_0 _26244_ (.A1(_07206_),
    .A2(_07459_),
    .B1(_07313_),
    .Y(_07460_));
 sky130_fd_sc_hd__inv_2 _26245_ (.A(_07194_),
    .Y(\if_stage_i.compressed_decoder_i.is_compressed_o ));
 sky130_fd_sc_hd__nor2_1 _26246_ (.A(_10842_),
    .B(\if_stage_i.compressed_decoder_i.is_compressed_o ),
    .Y(_07461_));
 sky130_fd_sc_hd__o21ai_0 _26247_ (.A1(_10867_),
    .A2(_07179_),
    .B1(_10842_),
    .Y(_07462_));
 sky130_fd_sc_hd__o21ai_0 _26248_ (.A1(_07190_),
    .A2(_07461_),
    .B1(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__nand2_2 _26249_ (.A(_07460_),
    .B(_07463_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[5] ));
 sky130_fd_sc_hd__nor2_1 _26250_ (.A(_10776_),
    .B(_07409_),
    .Y(_07464_));
 sky130_fd_sc_hd__a32oi_1 _26251_ (.A1(_07173_),
    .A2(_07163_),
    .A3(_07141_),
    .B1(_07464_),
    .B2(_10769_),
    .Y(_07465_));
 sky130_fd_sc_hd__o21ai_0 _26252_ (.A1(_10838_),
    .A2(_07437_),
    .B1(_07465_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[6] ));
 sky130_fd_sc_hd__nor2_1 _26253_ (.A(_10867_),
    .B(_10873_),
    .Y(_07466_));
 sky130_fd_sc_hd__o31ai_1 _26254_ (.A1(_10896_),
    .A2(_07155_),
    .A3(_07146_),
    .B1(_10879_),
    .Y(_07467_));
 sky130_fd_sc_hd__o21ai_0 _26255_ (.A1(_10878_),
    .A2(_07466_),
    .B1(\if_stage_i.compressed_decoder_i.instr_i[7] ),
    .Y(_07468_));
 sky130_fd_sc_hd__a21oi_1 _26256_ (.A1(_10898_),
    .A2(_07203_),
    .B1(_07368_),
    .Y(_07469_));
 sky130_fd_sc_hd__a21oi_1 _26257_ (.A1(_07468_),
    .A2(_07469_),
    .B1(_07137_),
    .Y(_07470_));
 sky130_fd_sc_hd__a31oi_1 _26258_ (.A1(_07163_),
    .A2(_07466_),
    .A3(_07467_),
    .B1(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__a21oi_1 _26259_ (.A1(_10776_),
    .A2(_07173_),
    .B1(_07140_),
    .Y(_07472_));
 sky130_fd_sc_hd__o21ai_0 _26260_ (.A1(_10867_),
    .A2(_07472_),
    .B1(_10767_),
    .Y(_07473_));
 sky130_fd_sc_hd__o21ai_0 _26261_ (.A1(_10769_),
    .A2(_07324_),
    .B1(_10776_),
    .Y(_07474_));
 sky130_fd_sc_hd__nand3_1 _26262_ (.A(_07471_),
    .B(_07473_),
    .C(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__o21ai_0 _26263_ (.A1(_07198_),
    .A2(_07471_),
    .B1(_10846_),
    .Y(_07476_));
 sky130_fd_sc_hd__a32o_1 _26264_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .A2(_07159_),
    .A3(_07151_),
    .B1(_07475_),
    .B2(_07476_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[7] ));
 sky130_fd_sc_hd__a21oi_1 _26265_ (.A1(_10872_),
    .A2(_07146_),
    .B1(_07287_),
    .Y(_07477_));
 sky130_fd_sc_hd__o22ai_1 _26266_ (.A1(_10767_),
    .A2(_07464_),
    .B1(_07477_),
    .B2(_10775_),
    .Y(_07478_));
 sky130_fd_sc_hd__a32oi_1 _26267_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .A2(_07203_),
    .A3(_07313_),
    .B1(_07478_),
    .B2(_10850_),
    .Y(_07479_));
 sky130_fd_sc_hd__a221oi_1 _26268_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .A2(_07159_),
    .B1(_07271_),
    .B2(_10850_),
    .C1(_07248_),
    .Y(_07480_));
 sky130_fd_sc_hd__a21oi_1 _26269_ (.A1(_07248_),
    .A2(_07479_),
    .B1(_07480_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[8] ));
 sky130_fd_sc_hd__a32oi_1 _26270_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .A2(_10866_),
    .A3(_07203_),
    .B1(_07271_),
    .B2(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .Y(_07481_));
 sky130_fd_sc_hd__o22ai_1 _26271_ (.A1(_07157_),
    .A2(_07248_),
    .B1(_07233_),
    .B2(_07137_),
    .Y(_07482_));
 sky130_fd_sc_hd__a32oi_1 _26272_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .A2(_07263_),
    .A3(_07409_),
    .B1(_07482_),
    .B2(_10892_),
    .Y(_07483_));
 sky130_fd_sc_hd__nand3_1 _26273_ (.A(_10776_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .C(_07174_),
    .Y(_07484_));
 sky130_fd_sc_hd__o211ai_1 _26274_ (.A1(_07248_),
    .A2(_07481_),
    .B1(_07483_),
    .C1(_07484_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[9] ));
 sky130_fd_sc_hd__inv_1 _26275_ (.A(net94),
    .Y(_07485_));
 sky130_fd_sc_hd__o21ai_0 _26276_ (.A1(_07485_),
    .A2(_10916_),
    .B1(_10908_),
    .Y(_07486_));
 sky130_fd_sc_hd__nand2_1 _26277_ (.A(net3948),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__a211oi_1 _26278_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(_10918_),
    .B1(_07066_),
    .C1(_10908_),
    .Y(_07488_));
 sky130_fd_sc_hd__a21oi_1 _26279_ (.A1(_10917_),
    .A2(_07487_),
    .B1(_07488_),
    .Y(\if_stage_i.fetch_err ));
 sky130_fd_sc_hd__a21oi_1 _26280_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(net3567),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .Y(_07489_));
 sky130_fd_sc_hd__o21ai_0 _26281_ (.A1(net128),
    .A2(net3567),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Y(_07490_));
 sky130_fd_sc_hd__inv_1 _26282_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .Y(_07491_));
 sky130_fd_sc_hd__a32oi_1 _26283_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .A3(_07489_),
    .B1(_07490_),
    .B2(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__a21o_1 _26284_ (.A1(net95),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .B1(_07492_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 sky130_fd_sc_hd__nand3_1 _26285_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(net95),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Y(_07493_));
 sky130_fd_sc_hd__a21boi_0 _26286_ (.A1(_07489_),
    .A2(_07493_),
    .B1_N(_10912_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 sky130_fd_sc_hd__a31oi_4 _26287_ (.A1(net3742),
    .A2(_10646_),
    .A3(_10781_),
    .B1(_10825_),
    .Y(_07494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__o21ai_0 _26290_ (.A1(_10642_),
    .A2(_10784_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Y(_07497_));
 sky130_fd_sc_hd__a21oi_1 _26291_ (.A1(_10495_),
    .A2(_07497_),
    .B1(_10538_),
    .Y(_07498_));
 sky130_fd_sc_hd__or2_4 _26292_ (.A(_12176_),
    .B(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__or2_4 _26293_ (.A(_12181_),
    .B(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_48 ();
 sky130_fd_sc_hd__nor2_1 _26295_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10784_),
    .Y(_07502_));
 sky130_fd_sc_hd__o21ai_4 _26296_ (.A1(_10782_),
    .A2(_07502_),
    .B1(_12171_),
    .Y(_07503_));
 sky130_fd_sc_hd__nand2_4 _26297_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_12754_),
    .Y(_07504_));
 sky130_fd_sc_hd__and3_4 _26298_ (.A(_12171_),
    .B(_07503_),
    .C(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__a222oi_1 _26300_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[10] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[10] ),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_1 _26301_ (.A(net3515),
    .B(net3742),
    .Y(_07508_));
 sky130_fd_sc_hd__nor2_1 _26302_ (.A(net1),
    .B(_07500_),
    .Y(_07509_));
 sky130_fd_sc_hd__a31oi_2 _26303_ (.A1(_07500_),
    .A2(_07507_),
    .A3(_07508_),
    .B1(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_1 _26304_ (.A(net3567),
    .B(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__a21boi_2 _26305_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .A2(net3554),
    .B1_N(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__inv_1 _26306_ (.A(\cs_registers_i.csr_depc_o[7] ),
    .Y(_07513_));
 sky130_fd_sc_hd__a21oi_1 _26307_ (.A1(_07513_),
    .A2(_12181_),
    .B1(_07499_),
    .Y(_07514_));
 sky130_fd_sc_hd__a221oi_2 _26308_ (.A1(net178),
    .A2(net3742),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .C1(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__nand2_2 _26309_ (.A(net3567),
    .B(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__o21ai_2 _26310_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .A2(net3567),
    .B1(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__a221oi_2 _26311_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[6] ),
    .C1(_12481_),
    .Y(_07518_));
 sky130_fd_sc_hd__o21ai_4 _26312_ (.A1(net3529),
    .A2(_10540_),
    .B1(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nor2_4 _26313_ (.A(_12181_),
    .B(_07499_),
    .Y(_07520_));
 sky130_fd_sc_hd__nor2_2 _26314_ (.A(net3554),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__a22oi_2 _26315_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(net3554),
    .B1(_07519_),
    .B2(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand2_4 _26316_ (.A(_10826_),
    .B(_07500_),
    .Y(_07523_));
 sky130_fd_sc_hd__a22oi_2 _26317_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .Y(_07524_));
 sky130_fd_sc_hd__nand2_2 _26318_ (.A(_12471_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__a21oi_4 _26319_ (.A1(net3742),
    .A2(net3537),
    .B1(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__nor2_2 _26320_ (.A(_07523_),
    .B(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__a21oi_2 _26321_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .A2(_07494_),
    .B1(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__a22oi_1 _26322_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .Y(_07529_));
 sky130_fd_sc_hd__nand2_1 _26323_ (.A(net3742),
    .B(net3535),
    .Y(_07530_));
 sky130_fd_sc_hd__nand4_1 _26324_ (.A(_10826_),
    .B(_12465_),
    .C(_07529_),
    .D(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__o21a_1 _26325_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .A2(net3567),
    .B1(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__inv_1 _26326_ (.A(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__a22oi_2 _26327_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(_12181_),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .Y(_07534_));
 sky130_fd_sc_hd__nand3_2 _26328_ (.A(_12450_),
    .B(_07504_),
    .C(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__a21oi_2 _26329_ (.A1(net3742),
    .A2(net174),
    .B1(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__nor2_2 _26330_ (.A(_07523_),
    .B(_07536_),
    .Y(_07537_));
 sky130_fd_sc_hd__a21oi_2 _26331_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .A2(_07494_),
    .B1(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__a221oi_4 _26332_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_12181_),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[2] ),
    .C1(_12433_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_2 _26333_ (.A(net3742),
    .B(net171),
    .Y(_07540_));
 sky130_fd_sc_hd__a21oi_4 _26334_ (.A1(_07539_),
    .A2(_07540_),
    .B1(_07523_),
    .Y(_07541_));
 sky130_fd_sc_hd__and2_4 _26335_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .B(_07494_),
    .X(_07542_));
 sky130_fd_sc_hd__nor2_2 _26336_ (.A(_07541_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__nand2b_4 _26337_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_07070_),
    .Y(_07544_));
 sky130_fd_sc_hd__or3_4 _26338_ (.A(_07538_),
    .B(_07543_),
    .C(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__or3_4 _26339_ (.A(_07528_),
    .B(_07533_),
    .C(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__or3_4 _26340_ (.A(_07517_),
    .B(_07522_),
    .C(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__nand2_1 _26342_ (.A(\cs_registers_i.csr_mtvec_o[9] ),
    .B(_07505_),
    .Y(_07549_));
 sky130_fd_sc_hd__a22oi_1 _26343_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .Y(_07550_));
 sky130_fd_sc_hd__nand2_2 _26344_ (.A(_07549_),
    .B(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__nand2_1 _26345_ (.A(\cs_registers_i.csr_mtvec_o[8] ),
    .B(_07505_),
    .Y(_07552_));
 sky130_fd_sc_hd__a22oi_1 _26346_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[8] ),
    .Y(_07553_));
 sky130_fd_sc_hd__nand2_2 _26347_ (.A(_07552_),
    .B(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__a21oi_1 _26348_ (.A1(_07551_),
    .A2(_07554_),
    .B1(net3742),
    .Y(_07555_));
 sky130_fd_sc_hd__o22ai_1 _26349_ (.A1(net3520),
    .A2(_07551_),
    .B1(_07554_),
    .B2(net3519),
    .Y(_07556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__nand3_1 _26351_ (.A(net23),
    .B(net24),
    .C(_07520_),
    .Y(_07558_));
 sky130_fd_sc_hd__o21ai_2 _26352_ (.A1(_07555_),
    .A2(_07556_),
    .B1(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__and3_1 _26353_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .C(net3554),
    .X(_07560_));
 sky130_fd_sc_hd__a21oi_2 _26354_ (.A1(net3567),
    .A2(_07559_),
    .B1(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__nor3_1 _26355_ (.A(_07512_),
    .B(_07547_),
    .C(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__o21a_1 _26356_ (.A1(_07547_),
    .A2(_07561_),
    .B1(_07512_),
    .X(_07563_));
 sky130_fd_sc_hd__nor2_1 _26357_ (.A(_07562_),
    .B(_07563_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ));
 sky130_fd_sc_hd__nor2_1 _26358_ (.A(net2),
    .B(_07500_),
    .Y(_07564_));
 sky130_fd_sc_hd__nand2_8 _26359_ (.A(_12171_),
    .B(_07504_),
    .Y(_07565_));
 sky130_fd_sc_hd__o21ai_0 _26360_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07566_));
 sky130_fd_sc_hd__a22oi_1 _26361_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_12181_),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[11] ),
    .Y(_07567_));
 sky130_fd_sc_hd__nand2_2 _26362_ (.A(_07566_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__a211oi_1 _26363_ (.A1(net3516),
    .A2(net3742),
    .B1(_07520_),
    .C1(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__nor3_2 _26364_ (.A(net3554),
    .B(_07564_),
    .C(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__a21oi_2 _26365_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .A2(net3554),
    .B1(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__xnor2_1 _26366_ (.A(_07562_),
    .B(_07571_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ));
 sky130_fd_sc_hd__nor4_1 _26367_ (.A(_07512_),
    .B(_07547_),
    .C(_07561_),
    .D(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__a222oi_1 _26368_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[12] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[12] ),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2_4 _26369_ (.A(net153),
    .B(net3742),
    .Y(_07574_));
 sky130_fd_sc_hd__nor2_1 _26370_ (.A(net3),
    .B(_07500_),
    .Y(_07575_));
 sky130_fd_sc_hd__a311oi_2 _26371_ (.A1(_07500_),
    .A2(_07573_),
    .A3(_07574_),
    .B1(_07575_),
    .C1(net3554),
    .Y(_07576_));
 sky130_fd_sc_hd__a21oi_2 _26372_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .A2(net3554),
    .B1(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__xnor2_1 _26373_ (.A(_07572_),
    .B(_07577_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ));
 sky130_fd_sc_hd__nand4_1 _26374_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .D(net3554),
    .Y(_07578_));
 sky130_fd_sc_hd__nand3_1 _26375_ (.A(net3567),
    .B(_07510_),
    .C(_07559_),
    .Y(_07579_));
 sky130_fd_sc_hd__a2111oi_0 _26376_ (.A1(_07578_),
    .A2(_07579_),
    .B1(_07577_),
    .C1(_07571_),
    .D1(_07547_),
    .Y(_07580_));
 sky130_fd_sc_hd__a222oi_1 _26377_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[13] ),
    .Y(_07581_));
 sky130_fd_sc_hd__nand2_1 _26378_ (.A(net4),
    .B(_07520_),
    .Y(_07582_));
 sky130_fd_sc_hd__o2111ai_4 _26379_ (.A1(net3498),
    .A2(_10540_),
    .B1(_10826_),
    .C1(_07581_),
    .D1(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__o21a_4 _26380_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .A2(net3567),
    .B1(_07583_),
    .X(_07584_));
 sky130_fd_sc_hd__xor2_1 _26381_ (.A(net3466),
    .B(_07584_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ));
 sky130_fd_sc_hd__nand2_8 _26382_ (.A(net155),
    .B(net3742),
    .Y(_07585_));
 sky130_fd_sc_hd__a222oi_1 _26383_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[14] ),
    .Y(_07586_));
 sky130_fd_sc_hd__nand2_1 _26384_ (.A(net5),
    .B(_07520_),
    .Y(_07587_));
 sky130_fd_sc_hd__nand4_1 _26385_ (.A(net3567),
    .B(_07585_),
    .C(_07586_),
    .D(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__o21a_4 _26386_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(net3567),
    .B1(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__and3b_4 _26387_ (.A_N(_07577_),
    .B(_07584_),
    .C(_07572_),
    .X(_07590_));
 sky130_fd_sc_hd__xor2_1 _26388_ (.A(_07589_),
    .B(_07590_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ));
 sky130_fd_sc_hd__a222oi_1 _26389_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(net3610),
    .B1(net3662),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[15] ),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _26390_ (.A(net6),
    .B(_07520_),
    .Y(_07592_));
 sky130_fd_sc_hd__nand3_1 _26391_ (.A(net3567),
    .B(_07591_),
    .C(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__a21oi_2 _26392_ (.A1(net3507),
    .A2(net3742),
    .B1(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nor2_1 _26393_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .B(net3567),
    .Y(_07595_));
 sky130_fd_sc_hd__nor2_1 _26394_ (.A(_07594_),
    .B(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__nand2_1 _26395_ (.A(_07589_),
    .B(_07590_),
    .Y(_07597_));
 sky130_fd_sc_hd__xnor2_1 _26396_ (.A(_07596_),
    .B(_07597_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ));
 sky130_fd_sc_hd__nand2_1 _26397_ (.A(net3506),
    .B(net3742),
    .Y(_07598_));
 sky130_fd_sc_hd__o21ai_0 _26398_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07599_));
 sky130_fd_sc_hd__a22oi_1 _26399_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[16] ),
    .Y(_07600_));
 sky130_fd_sc_hd__nand4_1 _26400_ (.A(_07500_),
    .B(_07598_),
    .C(_07599_),
    .D(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__o211ai_1 _26401_ (.A1(net7),
    .A2(_07500_),
    .B1(_07601_),
    .C1(_10826_),
    .Y(_07602_));
 sky130_fd_sc_hd__a21boi_4 _26402_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A2(net3554),
    .B1_N(net358),
    .Y(_07603_));
 sky130_fd_sc_hd__nand4_1 _26403_ (.A(net3466),
    .B(_07584_),
    .C(_07589_),
    .D(_07596_),
    .Y(_07604_));
 sky130_fd_sc_hd__xor2_1 _26404_ (.A(_07603_),
    .B(_07604_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ));
 sky130_fd_sc_hd__nor2_1 _26405_ (.A(_07603_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__nand2_2 _26406_ (.A(net158),
    .B(net3742),
    .Y(_07606_));
 sky130_fd_sc_hd__a222oi_1 _26407_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[17] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[17] ),
    .Y(_07607_));
 sky130_fd_sc_hd__nand2_1 _26408_ (.A(net8),
    .B(net3569),
    .Y(_07608_));
 sky130_fd_sc_hd__nand4_1 _26409_ (.A(_10826_),
    .B(_07606_),
    .C(_07607_),
    .D(_07608_),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_2 _26410_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(net3567),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__xnor2_1 _26411_ (.A(_07605_),
    .B(_07610_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__a222oi_1 _26413_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[18] ),
    .Y(_07612_));
 sky130_fd_sc_hd__nand2_1 _26414_ (.A(net9),
    .B(net3569),
    .Y(_07613_));
 sky130_fd_sc_hd__o2111ai_4 _26415_ (.A1(_10540_),
    .A2(net3497),
    .B1(_10826_),
    .C1(_07612_),
    .D1(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21ai_2 _26416_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .A2(net3567),
    .B1(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__nor3_1 _26417_ (.A(_07603_),
    .B(_07604_),
    .C(_07610_),
    .Y(_07616_));
 sky130_fd_sc_hd__xnor2_1 _26418_ (.A(_07615_),
    .B(_07616_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ));
 sky130_fd_sc_hd__nand2_4 _26419_ (.A(net160),
    .B(net3742),
    .Y(_07617_));
 sky130_fd_sc_hd__a222oi_1 _26420_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[19] ),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_1 _26421_ (.A(net10),
    .B(net3569),
    .Y(_07619_));
 sky130_fd_sc_hd__nand4_1 _26422_ (.A(_10826_),
    .B(_07617_),
    .C(_07618_),
    .D(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__o21a_4 _26423_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(net3567),
    .B1(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__nor4_2 _26424_ (.A(_07603_),
    .B(_07604_),
    .C(_07610_),
    .D(_07615_),
    .Y(_07622_));
 sky130_fd_sc_hd__xor2_1 _26425_ (.A(_07621_),
    .B(net3454),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ));
 sky130_fd_sc_hd__nand2_1 _26426_ (.A(net11),
    .B(net3569),
    .Y(_07623_));
 sky130_fd_sc_hd__o21ai_0 _26427_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07624_));
 sky130_fd_sc_hd__a22oi_1 _26428_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[20] ),
    .Y(_07625_));
 sky130_fd_sc_hd__nand4_1 _26429_ (.A(_10826_),
    .B(_07623_),
    .C(_07624_),
    .D(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a21oi_4 _26430_ (.A1(net3505),
    .A2(net3742),
    .B1(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__nor2_1 _26431_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .B(net3567),
    .Y(_07628_));
 sky130_fd_sc_hd__nor2_2 _26432_ (.A(_07627_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_1 _26433_ (.A(_07621_),
    .B(net3454),
    .Y(_07630_));
 sky130_fd_sc_hd__xnor2_1 _26434_ (.A(_07629_),
    .B(_07630_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ));
 sky130_fd_sc_hd__a222oi_1 _26435_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[21] ),
    .Y(_07631_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__nand2_1 _26437_ (.A(net12),
    .B(_07520_),
    .Y(_07633_));
 sky130_fd_sc_hd__o2111ai_2 _26438_ (.A1(net3496),
    .A2(_10540_),
    .B1(net3567),
    .C1(_07631_),
    .D1(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__o21a_1 _26439_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .A2(net3567),
    .B1(_07634_),
    .X(_07635_));
 sky130_fd_sc_hd__nand3_4 _26440_ (.A(_07621_),
    .B(_07622_),
    .C(_07629_),
    .Y(_07636_));
 sky130_fd_sc_hd__xnor2_1 _26441_ (.A(_07635_),
    .B(_07636_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ));
 sky130_fd_sc_hd__nand2_2 _26442_ (.A(net3503),
    .B(net3742),
    .Y(_07637_));
 sky130_fd_sc_hd__a222oi_1 _26443_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[22] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[22] ),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _26444_ (.A(net13),
    .B(net3569),
    .Y(_07639_));
 sky130_fd_sc_hd__nand4_1 _26445_ (.A(_10826_),
    .B(_07637_),
    .C(_07638_),
    .D(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__o21a_4 _26446_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(net3567),
    .B1(net377),
    .X(_07641_));
 sky130_fd_sc_hd__o21ai_1 _26447_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .A2(net3567),
    .B1(_07634_),
    .Y(_07642_));
 sky130_fd_sc_hd__nor2_1 _26448_ (.A(_07642_),
    .B(_07636_),
    .Y(_07643_));
 sky130_fd_sc_hd__xor2_1 _26449_ (.A(_07641_),
    .B(_07643_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ));
 sky130_fd_sc_hd__a222oi_1 _26450_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[23] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[23] ),
    .Y(_07644_));
 sky130_fd_sc_hd__nand2_1 _26451_ (.A(net14),
    .B(net3569),
    .Y(_07645_));
 sky130_fd_sc_hd__o2111ai_4 _26452_ (.A1(net3504),
    .A2(_10540_),
    .B1(_10826_),
    .C1(_07644_),
    .D1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__o21ai_2 _26453_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .A2(net3567),
    .B1(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__nand2_1 _26454_ (.A(_07635_),
    .B(_07641_),
    .Y(_07648_));
 sky130_fd_sc_hd__nor2_1 _26455_ (.A(_07636_),
    .B(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__xnor2_1 _26456_ (.A(_07647_),
    .B(_07649_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ));
 sky130_fd_sc_hd__nand2_2 _26457_ (.A(net273),
    .B(net3742),
    .Y(_07650_));
 sky130_fd_sc_hd__a222oi_1 _26458_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[24] ),
    .Y(_07651_));
 sky130_fd_sc_hd__nand2_1 _26459_ (.A(net15),
    .B(_07520_),
    .Y(_07652_));
 sky130_fd_sc_hd__nand4_1 _26460_ (.A(net3567),
    .B(_07650_),
    .C(_07651_),
    .D(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__o21ai_2 _26461_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(net3567),
    .B1(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__nor3_1 _26462_ (.A(_07636_),
    .B(_07647_),
    .C(_07648_),
    .Y(_07655_));
 sky130_fd_sc_hd__xnor2_1 _26463_ (.A(_07654_),
    .B(_07655_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ));
 sky130_fd_sc_hd__o21ai_0 _26464_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07656_));
 sky130_fd_sc_hd__a22oi_1 _26465_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .Y(_07657_));
 sky130_fd_sc_hd__nand2_1 _26466_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_2 _26467_ (.A1(net16),
    .A2(net3569),
    .B1(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__nand2_4 _26468_ (.A(net3495),
    .B(net3742),
    .Y(_07660_));
 sky130_fd_sc_hd__nand3_4 _26469_ (.A(_10826_),
    .B(_07659_),
    .C(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__o21a_4 _26470_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .A2(net3567),
    .B1(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__nor4_1 _26471_ (.A(_07636_),
    .B(_07647_),
    .C(_07648_),
    .D(_07654_),
    .Y(_07663_));
 sky130_fd_sc_hd__xor2_1 _26472_ (.A(_07662_),
    .B(_07663_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ));
 sky130_fd_sc_hd__a222oi_1 _26473_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[26] ),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_2 _26474_ (.A(net17),
    .B(_07520_),
    .Y(_07665_));
 sky130_fd_sc_hd__o2111ai_4 _26475_ (.A1(net3486),
    .A2(_10540_),
    .B1(net3567),
    .C1(_07664_),
    .D1(_07665_),
    .Y(_07666_));
 sky130_fd_sc_hd__o21a_4 _26476_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(net3567),
    .B1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__and2_4 _26477_ (.A(_07662_),
    .B(_07663_),
    .X(_07668_));
 sky130_fd_sc_hd__xor2_1 _26478_ (.A(_07667_),
    .B(_07668_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ));
 sky130_fd_sc_hd__o21ai_0 _26479_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07669_));
 sky130_fd_sc_hd__a22oi_1 _26480_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .Y(_07670_));
 sky130_fd_sc_hd__nand2_1 _26481_ (.A(_07669_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__a211oi_1 _26482_ (.A1(net18),
    .A2(_07520_),
    .B1(_07671_),
    .C1(net3554),
    .Y(_07672_));
 sky130_fd_sc_hd__o21ai_2 _26483_ (.A1(net3487),
    .A2(_10540_),
    .B1(_07672_),
    .Y(_07673_));
 sky130_fd_sc_hd__o21a_4 _26484_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .A2(net3567),
    .B1(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__nand2_1 _26485_ (.A(_07667_),
    .B(_07668_),
    .Y(_07675_));
 sky130_fd_sc_hd__xnor2_1 _26486_ (.A(_07674_),
    .B(_07675_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ));
 sky130_fd_sc_hd__nand2_1 _26487_ (.A(net19),
    .B(_07520_),
    .Y(_07676_));
 sky130_fd_sc_hd__o21ai_0 _26488_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_07565_),
    .B1(_07503_),
    .Y(_07677_));
 sky130_fd_sc_hd__a22oi_1 _26489_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .Y(_07678_));
 sky130_fd_sc_hd__nand4_1 _26490_ (.A(net3567),
    .B(_07676_),
    .C(_07677_),
    .D(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__a21oi_4 _26491_ (.A1(net169),
    .A2(net3742),
    .B1(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__o21bai_2 _26492_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .A2(net3567),
    .B1_N(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__nand3_1 _26493_ (.A(_07667_),
    .B(_07668_),
    .C(_07674_),
    .Y(_07682_));
 sky130_fd_sc_hd__xor2_1 _26494_ (.A(_07681_),
    .B(_07682_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ));
 sky130_fd_sc_hd__nand2_8 _26495_ (.A(net3742),
    .B(net170),
    .Y(_07683_));
 sky130_fd_sc_hd__a222oi_1 _26496_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(net3610),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[29] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[29] ),
    .Y(_07684_));
 sky130_fd_sc_hd__nand2_1 _26497_ (.A(net20),
    .B(_07520_),
    .Y(_07685_));
 sky130_fd_sc_hd__nand4_1 _26498_ (.A(net3567),
    .B(_07685_),
    .C(_07684_),
    .D(_07683_),
    .Y(_07686_));
 sky130_fd_sc_hd__o21ai_2 _26499_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .A2(net3567),
    .B1(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__or2_4 _26500_ (.A(_07681_),
    .B(_07682_),
    .X(_07688_));
 sky130_fd_sc_hd__xor2_1 _26501_ (.A(net466),
    .B(_07688_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ));
 sky130_fd_sc_hd__xor2_1 _26502_ (.A(_07543_),
    .B(_07544_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 sky130_fd_sc_hd__nand2_4 _26503_ (.A(net3473),
    .B(net3742),
    .Y(_07689_));
 sky130_fd_sc_hd__a222oi_1 _26504_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(net3611),
    .B1(net3663),
    .B2(\cs_registers_i.csr_mepc_o[30] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[30] ),
    .Y(_07690_));
 sky130_fd_sc_hd__nand2_1 _26505_ (.A(net21),
    .B(net3569),
    .Y(_07691_));
 sky130_fd_sc_hd__nand4_1 _26506_ (.A(_10826_),
    .B(_07689_),
    .C(_07690_),
    .D(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__o21a_4 _26507_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .A2(net3567),
    .B1(net271),
    .X(_07693_));
 sky130_fd_sc_hd__nor2_1 _26508_ (.A(net466),
    .B(_07688_),
    .Y(_07694_));
 sky130_fd_sc_hd__xor2_1 _26509_ (.A(_07693_),
    .B(_07694_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ));
 sky130_fd_sc_hd__a222oi_1 _26510_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[31] ),
    .C1(_07505_),
    .C2(\cs_registers_i.csr_mtvec_o[31] ),
    .Y(_07695_));
 sky130_fd_sc_hd__nand2_1 _26511_ (.A(net22),
    .B(net3569),
    .Y(_07696_));
 sky130_fd_sc_hd__o2111ai_4 _26512_ (.A1(net3471),
    .A2(_10540_),
    .B1(_10826_),
    .C1(_07695_),
    .D1(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__o21ai_4 _26513_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .A2(net3567),
    .B1(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand2_1 _26514_ (.A(_07693_),
    .B(_07694_),
    .Y(_07699_));
 sky130_fd_sc_hd__xor2_1 _26515_ (.A(_07698_),
    .B(_07699_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ));
 sky130_fd_sc_hd__o21ai_0 _26516_ (.A1(_07543_),
    .A2(_07544_),
    .B1(_07538_),
    .Y(_07700_));
 sky130_fd_sc_hd__and2_0 _26517_ (.A(_07545_),
    .B(_07700_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 sky130_fd_sc_hd__xnor2_1 _26518_ (.A(_07532_),
    .B(_07545_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ));
 sky130_fd_sc_hd__o21ai_0 _26519_ (.A1(_07533_),
    .A2(_07545_),
    .B1(_07528_),
    .Y(_07701_));
 sky130_fd_sc_hd__and2_0 _26520_ (.A(_07546_),
    .B(_07701_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ));
 sky130_fd_sc_hd__xor2_1 _26521_ (.A(_07522_),
    .B(_07546_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ));
 sky130_fd_sc_hd__nor2_1 _26522_ (.A(_07522_),
    .B(_07546_),
    .Y(_07702_));
 sky130_fd_sc_hd__xnor2_1 _26523_ (.A(_07517_),
    .B(_07702_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ));
 sky130_fd_sc_hd__a21oi_1 _26524_ (.A1(net3519),
    .A2(net3742),
    .B1(_07554_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_1 _26525_ (.A(_07500_),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__o21ai_2 _26526_ (.A1(net23),
    .A2(_07500_),
    .B1(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__nor2_2 _26527_ (.A(net3554),
    .B(_07705_),
    .Y(_07706_));
 sky130_fd_sc_hd__a21oi_2 _26528_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(net3554),
    .B1(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__xor2_1 _26529_ (.A(_07547_),
    .B(_07707_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__inv_1 _26531_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .Y(_07709_));
 sky130_fd_sc_hd__nor2_1 _26532_ (.A(_07709_),
    .B(_07547_),
    .Y(_07710_));
 sky130_fd_sc_hd__xnor2_1 _26533_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__a21oi_1 _26534_ (.A1(net3520),
    .A2(net3742),
    .B1(_07551_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand2_1 _26535_ (.A(_07500_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__o21ai_2 _26536_ (.A1(net24),
    .A2(_07500_),
    .B1(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__nor2_1 _26537_ (.A(_07547_),
    .B(_07705_),
    .Y(_07715_));
 sky130_fd_sc_hd__xnor2_1 _26538_ (.A(_07714_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand2_1 _26539_ (.A(net3567),
    .B(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__o21ai_0 _26540_ (.A1(net3567),
    .A2(_07711_),
    .B1(_07717_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__nand2_8 _26542_ (.A(net3554),
    .B(_07544_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ));
 sky130_fd_sc_hd__a21oi_1 _26543_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .Y(_07719_));
 sky130_fd_sc_hd__a211oi_1 _26544_ (.A1(net107),
    .A2(net96),
    .B1(net94),
    .C1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_07720_));
 sky130_fd_sc_hd__a21oi_2 _26545_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .A2(_07719_),
    .B1(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__nor2_4 _26546_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__nor2b_4 _26547_ (.A(_07722_),
    .B_N(_00009_),
    .Y(_07723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__nand2_1 _26549_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(_07723_),
    .Y(_07725_));
 sky130_fd_sc_hd__xnor2_1 _26550_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_07723_),
    .Y(_07726_));
 sky130_fd_sc_hd__nand2_4 _26551_ (.A(_10914_),
    .B(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__nand2_8 _26552_ (.A(net3414),
    .B(_07727_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ));
 sky130_fd_sc_hd__nand2b_1 _26553_ (.A_N(_07723_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_07728_));
 sky130_fd_sc_hd__o21ai_0 _26554_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_07728_),
    .B1(_07725_),
    .Y(_07729_));
 sky130_fd_sc_hd__a22o_4 _26555_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net3421),
    .B1(_07729_),
    .B2(_10914_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ));
 sky130_fd_sc_hd__o21ai_0 _26556_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_07485_),
    .B1(_07064_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ));
 sky130_fd_sc_hd__nand2_1 _26557_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .Y(_07730_));
 sky130_fd_sc_hd__o21ai_0 _26558_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(_07485_),
    .B1(_07730_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ));
 sky130_fd_sc_hd__a222oi_1 _26559_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(net3611),
    .B1(_12396_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .C1(_06418_),
    .C2(net3742),
    .Y(_07731_));
 sky130_fd_sc_hd__nor3b_1 _26560_ (.A(_07722_),
    .B(net3567),
    .C_N(_10919_),
    .Y(_07732_));
 sky130_fd_sc_hd__a21oi_1 _26561_ (.A1(net3567),
    .A2(_07731_),
    .B1(_07732_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[0] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__inv_1 _26563_ (.A(\cs_registers_i.pc_if_i[9] ),
    .Y(_07734_));
 sky130_fd_sc_hd__nand2_1 _26564_ (.A(\cs_registers_i.pc_if_i[5] ),
    .B(\cs_registers_i.pc_if_i[6] ),
    .Y(_07735_));
 sky130_fd_sc_hd__nor2b_4 _26565_ (.A(_07722_),
    .B_N(\cs_registers_i.pc_if_i[2] ),
    .Y(_07736_));
 sky130_fd_sc_hd__nand3_2 _26566_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__nor2_2 _26567_ (.A(_07735_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand3_2 _26568_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(\cs_registers_i.pc_if_i[8] ),
    .C(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__nor2_2 _26569_ (.A(_07734_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _26570_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__xnor2_1 _26571_ (.A(\cs_registers_i.pc_if_i[11] ),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__a21o_1 _26572_ (.A1(net3554),
    .A2(_07742_),
    .B1(_07570_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ));
 sky130_fd_sc_hd__nand3_2 _26573_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(\cs_registers_i.pc_if_i[11] ),
    .C(_07740_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_1 _26574_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__a21o_1 _26575_ (.A1(net3554),
    .A2(_07744_),
    .B1(_07576_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ));
 sky130_fd_sc_hd__inv_1 _26576_ (.A(\cs_registers_i.pc_if_i[12] ),
    .Y(_07745_));
 sky130_fd_sc_hd__nor2_2 _26577_ (.A(_07745_),
    .B(_07743_),
    .Y(_07746_));
 sky130_fd_sc_hd__xnor2_1 _26578_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__a21boi_0 _26579_ (.A1(net3554),
    .A2(_07747_),
    .B1_N(_07583_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ));
 sky130_fd_sc_hd__nand2_1 _26580_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_07746_),
    .Y(_07748_));
 sky130_fd_sc_hd__xor2_1 _26581_ (.A(\cs_registers_i.pc_if_i[14] ),
    .B(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__a21boi_0 _26582_ (.A1(net3554),
    .A2(_07749_),
    .B1_N(_07588_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ));
 sky130_fd_sc_hd__clkinv_1 _26583_ (.A(\cs_registers_i.pc_if_i[15] ),
    .Y(_07750_));
 sky130_fd_sc_hd__nand3_2 _26584_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(\cs_registers_i.pc_if_i[14] ),
    .C(_07746_),
    .Y(_07751_));
 sky130_fd_sc_hd__xnor2_1 _26585_ (.A(_07750_),
    .B(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__a21oi_1 _26586_ (.A1(net3554),
    .A2(_07752_),
    .B1(_07594_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ));
 sky130_fd_sc_hd__nor2_2 _26587_ (.A(_07750_),
    .B(_07751_),
    .Y(_07753_));
 sky130_fd_sc_hd__xnor2_1 _26588_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B(_07753_),
    .Y(_07754_));
 sky130_fd_sc_hd__o21ai_0 _26589_ (.A1(net3567),
    .A2(_07754_),
    .B1(net358),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ));
 sky130_fd_sc_hd__nand2_1 _26590_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B(_07753_),
    .Y(_07755_));
 sky130_fd_sc_hd__xor2_1 _26591_ (.A(\cs_registers_i.pc_if_i[17] ),
    .B(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__a21boi_0 _26592_ (.A1(net3554),
    .A2(_07756_),
    .B1_N(_07609_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ));
 sky130_fd_sc_hd__clkinv_1 _26593_ (.A(\cs_registers_i.pc_if_i[18] ),
    .Y(_07757_));
 sky130_fd_sc_hd__nand3_2 _26594_ (.A(\cs_registers_i.pc_if_i[16] ),
    .B(\cs_registers_i.pc_if_i[17] ),
    .C(_07753_),
    .Y(_07758_));
 sky130_fd_sc_hd__xnor2_1 _26595_ (.A(_07757_),
    .B(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__a21boi_0 _26596_ (.A1(net3554),
    .A2(_07759_),
    .B1_N(_07614_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__nor2_2 _26598_ (.A(_07757_),
    .B(_07758_),
    .Y(_07761_));
 sky130_fd_sc_hd__xnor2_1 _26599_ (.A(\cs_registers_i.pc_if_i[19] ),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__a21boi_0 _26600_ (.A1(net3554),
    .A2(_07762_),
    .B1_N(_07620_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ));
 sky130_fd_sc_hd__nand2_1 _26601_ (.A(\cs_registers_i.pc_if_i[19] ),
    .B(_07761_),
    .Y(_07763_));
 sky130_fd_sc_hd__xor2_1 _26602_ (.A(\cs_registers_i.pc_if_i[20] ),
    .B(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__a21oi_1 _26603_ (.A1(net3554),
    .A2(_07764_),
    .B1(_07627_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ));
 sky130_fd_sc_hd__xnor2_1 _26604_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_07722_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21o_1 _26605_ (.A1(net3554),
    .A2(_07765_),
    .B1(_07541_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ));
 sky130_fd_sc_hd__clkinv_1 _26606_ (.A(\cs_registers_i.pc_if_i[21] ),
    .Y(_07766_));
 sky130_fd_sc_hd__nand3_2 _26607_ (.A(\cs_registers_i.pc_if_i[19] ),
    .B(\cs_registers_i.pc_if_i[20] ),
    .C(_07761_),
    .Y(_07767_));
 sky130_fd_sc_hd__xnor2_1 _26608_ (.A(_07766_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__a21boi_0 _26609_ (.A1(net3554),
    .A2(_07768_),
    .B1_N(_07634_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ));
 sky130_fd_sc_hd__nor2_2 _26610_ (.A(_07766_),
    .B(_07767_),
    .Y(_07769_));
 sky130_fd_sc_hd__xnor2_1 _26611_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__a21boi_0 _26612_ (.A1(net3554),
    .A2(_07770_),
    .B1_N(net377),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ));
 sky130_fd_sc_hd__nand2_1 _26613_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B(_07769_),
    .Y(_07771_));
 sky130_fd_sc_hd__xor2_1 _26614_ (.A(\cs_registers_i.pc_if_i[23] ),
    .B(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__a21boi_0 _26615_ (.A1(net3554),
    .A2(_07772_),
    .B1_N(_07646_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ));
 sky130_fd_sc_hd__clkinv_1 _26616_ (.A(\cs_registers_i.pc_if_i[24] ),
    .Y(_07773_));
 sky130_fd_sc_hd__nand3_2 _26617_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B(\cs_registers_i.pc_if_i[23] ),
    .C(_07769_),
    .Y(_07774_));
 sky130_fd_sc_hd__xnor2_1 _26618_ (.A(_07773_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__a21boi_0 _26619_ (.A1(net3554),
    .A2(_07775_),
    .B1_N(_07653_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ));
 sky130_fd_sc_hd__nor2_2 _26620_ (.A(_07773_),
    .B(_07774_),
    .Y(_07776_));
 sky130_fd_sc_hd__xnor2_1 _26621_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__a21boi_0 _26622_ (.A1(net3554),
    .A2(_07777_),
    .B1_N(_07661_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ));
 sky130_fd_sc_hd__nand2_1 _26623_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B(_07776_),
    .Y(_07778_));
 sky130_fd_sc_hd__xor2_1 _26624_ (.A(\cs_registers_i.pc_if_i[26] ),
    .B(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__a21boi_0 _26625_ (.A1(net3554),
    .A2(_07779_),
    .B1_N(_07666_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ));
 sky130_fd_sc_hd__and3_4 _26626_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B(\cs_registers_i.pc_if_i[26] ),
    .C(_07776_),
    .X(_07780_));
 sky130_fd_sc_hd__xnor2_1 _26627_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__a21boi_0 _26628_ (.A1(net3554),
    .A2(_07781_),
    .B1_N(_07673_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ));
 sky130_fd_sc_hd__and2_4 _26629_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B(_07780_),
    .X(_07782_));
 sky130_fd_sc_hd__xnor2_1 _26630_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__a21oi_1 _26631_ (.A1(net3554),
    .A2(_07783_),
    .B1(_07680_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ));
 sky130_fd_sc_hd__nand2_1 _26632_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(_07782_),
    .Y(_07784_));
 sky130_fd_sc_hd__xor2_1 _26633_ (.A(\cs_registers_i.pc_if_i[29] ),
    .B(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__a21boi_0 _26634_ (.A1(net3554),
    .A2(_07785_),
    .B1_N(net441),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ));
 sky130_fd_sc_hd__nand3_1 _26635_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(\cs_registers_i.pc_if_i[29] ),
    .C(_07782_),
    .Y(_07786_));
 sky130_fd_sc_hd__xor2_1 _26636_ (.A(\cs_registers_i.pc_if_i[30] ),
    .B(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__a21boi_0 _26637_ (.A1(net3554),
    .A2(_07787_),
    .B1_N(net271),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ));
 sky130_fd_sc_hd__xnor2_1 _26638_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(_07736_),
    .Y(_07788_));
 sky130_fd_sc_hd__o22ai_1 _26639_ (.A1(_07523_),
    .A2(_07536_),
    .B1(_07788_),
    .B2(net3567),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ));
 sky130_fd_sc_hd__nand4_1 _26640_ (.A(\cs_registers_i.pc_if_i[28] ),
    .B(\cs_registers_i.pc_if_i[29] ),
    .C(\cs_registers_i.pc_if_i[30] ),
    .D(_07782_),
    .Y(_07789_));
 sky130_fd_sc_hd__xor2_1 _26641_ (.A(\cs_registers_i.pc_if_i[31] ),
    .B(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__a21boi_0 _26642_ (.A1(net3554),
    .A2(_07790_),
    .B1_N(_07697_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ));
 sky130_fd_sc_hd__a21o_1 _26643_ (.A1(\cs_registers_i.pc_if_i[3] ),
    .A2(_07736_),
    .B1(\cs_registers_i.pc_if_i[4] ),
    .X(_07791_));
 sky130_fd_sc_hd__nand2_1 _26644_ (.A(_07737_),
    .B(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__a21boi_0 _26645_ (.A1(net3554),
    .A2(_07792_),
    .B1_N(_07531_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ));
 sky130_fd_sc_hd__xor2_1 _26646_ (.A(\cs_registers_i.pc_if_i[5] ),
    .B(_07737_),
    .X(_07793_));
 sky130_fd_sc_hd__o22ai_1 _26647_ (.A1(_07523_),
    .A2(_07526_),
    .B1(_07793_),
    .B2(net3567),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ));
 sky130_fd_sc_hd__nand4_1 _26648_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(\cs_registers_i.pc_if_i[5] ),
    .D(_07736_),
    .Y(_07794_));
 sky130_fd_sc_hd__xor2_1 _26649_ (.A(\cs_registers_i.pc_if_i[6] ),
    .B(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__nand2_1 _26650_ (.A(_07519_),
    .B(_07521_),
    .Y(_07796_));
 sky130_fd_sc_hd__o21ai_0 _26651_ (.A1(net3567),
    .A2(_07795_),
    .B1(_07796_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ));
 sky130_fd_sc_hd__xnor2_1 _26652_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(_07738_),
    .Y(_07797_));
 sky130_fd_sc_hd__a21boi_0 _26653_ (.A1(net3554),
    .A2(_07797_),
    .B1_N(_07516_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ));
 sky130_fd_sc_hd__nand2_1 _26654_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(_07738_),
    .Y(_07798_));
 sky130_fd_sc_hd__xnor2_1 _26655_ (.A(\cs_registers_i.pc_if_i[8] ),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__a21o_1 _26656_ (.A1(net3554),
    .A2(_07799_),
    .B1(_07706_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ));
 sky130_fd_sc_hd__xnor2_1 _26657_ (.A(\cs_registers_i.pc_if_i[9] ),
    .B(_07739_),
    .Y(_07800_));
 sky130_fd_sc_hd__nor2_1 _26658_ (.A(net3554),
    .B(_07714_),
    .Y(_07801_));
 sky130_fd_sc_hd__a21o_1 _26659_ (.A1(net3554),
    .A2(_07800_),
    .B1(_07801_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ));
 sky130_fd_sc_hd__xnor2_1 _26660_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(_07740_),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ai_0 _26661_ (.A1(net3567),
    .A2(_07802_),
    .B1(_07511_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ));
 sky130_fd_sc_hd__nand2b_4 _26662_ (.A_N(net3440),
    .B(net3554),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ));
 sky130_fd_sc_hd__mux2_1 _26663_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ));
 sky130_fd_sc_hd__mux2_1 _26664_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ));
 sky130_fd_sc_hd__mux2_1 _26665_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ));
 sky130_fd_sc_hd__mux2_1 _26666_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ));
 sky130_fd_sc_hd__mux2_1 _26667_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ));
 sky130_fd_sc_hd__mux2_1 _26668_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__mux2_1 _26670_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ));
 sky130_fd_sc_hd__mux2_1 _26671_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ));
 sky130_fd_sc_hd__mux2_1 _26672_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ));
 sky130_fd_sc_hd__mux2_1 _26673_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ));
 sky130_fd_sc_hd__mux2_1 _26674_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ));
 sky130_fd_sc_hd__mux2_1 _26675_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ));
 sky130_fd_sc_hd__mux2_1 _26676_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ));
 sky130_fd_sc_hd__mux2_1 _26677_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ));
 sky130_fd_sc_hd__mux2_1 _26678_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ));
 sky130_fd_sc_hd__mux2_1 _26679_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ));
 sky130_fd_sc_hd__mux2_1 _26680_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ));
 sky130_fd_sc_hd__mux2_1 _26681_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ));
 sky130_fd_sc_hd__mux2_1 _26682_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ));
 sky130_fd_sc_hd__mux2_1 _26683_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__mux2_1 _26685_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ));
 sky130_fd_sc_hd__mux2_1 _26686_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ));
 sky130_fd_sc_hd__mux2_1 _26687_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ));
 sky130_fd_sc_hd__mux2_1 _26688_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ));
 sky130_fd_sc_hd__mux2_1 _26689_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ));
 sky130_fd_sc_hd__mux2_1 _26690_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ));
 sky130_fd_sc_hd__mux2_1 _26691_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ));
 sky130_fd_sc_hd__mux2_1 _26692_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ));
 sky130_fd_sc_hd__mux2_1 _26693_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ));
 sky130_fd_sc_hd__mux2_1 _26694_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__mux2_1 _26696_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ));
 sky130_fd_sc_hd__mux2_1 _26697_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ));
 sky130_fd_sc_hd__mux2_1 _26698_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ));
 sky130_fd_sc_hd__mux2_1 _26699_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ));
 sky130_fd_sc_hd__mux2_1 _26700_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ));
 sky130_fd_sc_hd__mux2_1 _26701_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ));
 sky130_fd_sc_hd__mux2_1 _26702_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ));
 sky130_fd_sc_hd__mux2_1 _26703_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ));
 sky130_fd_sc_hd__mux2_1 _26704_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ));
 sky130_fd_sc_hd__mux2_1 _26705_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ));
 sky130_fd_sc_hd__mux2_1 _26706_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ));
 sky130_fd_sc_hd__mux2_1 _26707_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ));
 sky130_fd_sc_hd__mux2_1 _26708_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ));
 sky130_fd_sc_hd__mux2_1 _26709_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ));
 sky130_fd_sc_hd__mux2_1 _26710_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ));
 sky130_fd_sc_hd__mux2_1 _26711_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ));
 sky130_fd_sc_hd__mux2_1 _26712_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ));
 sky130_fd_sc_hd__mux2_1 _26713_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ));
 sky130_fd_sc_hd__inv_1 _26714_ (.A(net3420),
    .Y(_07806_));
 sky130_fd_sc_hd__o311ai_0 _26715_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_10912_),
    .A3(net3420),
    .B1(net3414),
    .C1(_10913_),
    .Y(_07807_));
 sky130_fd_sc_hd__o311a_1 _26716_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_10914_),
    .A3(_07806_),
    .B1(_07807_),
    .C1(net3554),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 sky130_fd_sc_hd__nand2_1 _26717_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .B(net3419),
    .Y(_07808_));
 sky130_fd_sc_hd__nand3_1 _26718_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_10914_),
    .C(_07806_),
    .Y(_07809_));
 sky130_fd_sc_hd__o21ai_0 _26719_ (.A1(_10914_),
    .A2(_07806_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_07810_));
 sky130_fd_sc_hd__a31oi_1 _26720_ (.A1(_07808_),
    .A2(_07809_),
    .A3(_07810_),
    .B1(net3567),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 sky130_fd_sc_hd__a21oi_1 _26721_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_10914_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Y(_07811_));
 sky130_fd_sc_hd__nor3_1 _26722_ (.A(net3567),
    .B(net3419),
    .C(_07811_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 sky130_fd_sc_hd__inv_1 _26723_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .Y(_07812_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__mux2i_1 _26725_ (.A0(_07512_),
    .A1(_07812_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net219));
 sky130_fd_sc_hd__inv_1 _26726_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .Y(_07814_));
 sky130_fd_sc_hd__mux2i_1 _26727_ (.A0(_07571_),
    .A1(_07814_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net220));
 sky130_fd_sc_hd__inv_1 _26728_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .Y(_07815_));
 sky130_fd_sc_hd__mux2i_1 _26729_ (.A0(_07577_),
    .A1(_07815_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net221));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__mux2_1 _26731_ (.A0(_07584_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net222));
 sky130_fd_sc_hd__mux2_1 _26732_ (.A0(_07589_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net223));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__nand2_1 _26734_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .Y(_07818_));
 sky130_fd_sc_hd__o31ai_1 _26735_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07594_),
    .A3(_07595_),
    .B1(_07818_),
    .Y(net224));
 sky130_fd_sc_hd__inv_1 _26736_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .Y(_07819_));
 sky130_fd_sc_hd__mux2i_1 _26737_ (.A0(_07603_),
    .A1(_07819_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net225));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__nand2_1 _26739_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .Y(_07821_));
 sky130_fd_sc_hd__o21ai_0 _26740_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07610_),
    .B1(_07821_),
    .Y(net226));
 sky130_fd_sc_hd__nand2_1 _26741_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .Y(_07822_));
 sky130_fd_sc_hd__o21ai_1 _26742_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07615_),
    .B1(_07822_),
    .Y(net227));
 sky130_fd_sc_hd__mux2_1 _26743_ (.A0(_07621_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net228));
 sky130_fd_sc_hd__nand2_1 _26744_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .Y(_07823_));
 sky130_fd_sc_hd__o31ai_1 _26745_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07627_),
    .A3(_07628_),
    .B1(_07823_),
    .Y(net229));
 sky130_fd_sc_hd__nand2_1 _26746_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .Y(_07824_));
 sky130_fd_sc_hd__o21ai_0 _26747_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07642_),
    .B1(_07824_),
    .Y(net230));
 sky130_fd_sc_hd__mux2_1 _26748_ (.A0(_07641_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net231));
 sky130_fd_sc_hd__nand2_1 _26749_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .Y(_07825_));
 sky130_fd_sc_hd__o21ai_0 _26750_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07647_),
    .B1(_07825_),
    .Y(net232));
 sky130_fd_sc_hd__nand2_1 _26751_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .Y(_07826_));
 sky130_fd_sc_hd__o21ai_0 _26752_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07654_),
    .B1(_07826_),
    .Y(net233));
 sky130_fd_sc_hd__mux2_1 _26753_ (.A0(_07662_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net234));
 sky130_fd_sc_hd__mux2_1 _26754_ (.A0(_07667_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net235));
 sky130_fd_sc_hd__mux2_1 _26755_ (.A0(_07674_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net236));
 sky130_fd_sc_hd__nand2_1 _26756_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .Y(_07827_));
 sky130_fd_sc_hd__o21ai_0 _26757_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07681_),
    .B1(_07827_),
    .Y(net237));
 sky130_fd_sc_hd__nand2_1 _26758_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .Y(_07828_));
 sky130_fd_sc_hd__o21ai_2 _26759_ (.A1(_07687_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07828_),
    .Y(net238));
 sky130_fd_sc_hd__inv_1 _26760_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .Y(_07829_));
 sky130_fd_sc_hd__nor3_1 _26761_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_07541_),
    .C(_07542_),
    .Y(_07830_));
 sky130_fd_sc_hd__a21oi_1 _26762_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07829_),
    .B1(_07830_),
    .Y(net239));
 sky130_fd_sc_hd__mux2_2 _26763_ (.A0(_07693_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(net240));
 sky130_fd_sc_hd__nand2_1 _26764_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .Y(_07831_));
 sky130_fd_sc_hd__o21ai_2 _26765_ (.A1(_07698_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07831_),
    .Y(net241));
 sky130_fd_sc_hd__inv_1 _26766_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .Y(_07832_));
 sky130_fd_sc_hd__mux2i_1 _26767_ (.A0(_07538_),
    .A1(_07832_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net242));
 sky130_fd_sc_hd__nand2_1 _26768_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .Y(_07833_));
 sky130_fd_sc_hd__o21ai_0 _26769_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07533_),
    .B1(_07833_),
    .Y(net243));
 sky130_fd_sc_hd__inv_1 _26770_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .Y(_07834_));
 sky130_fd_sc_hd__mux2i_1 _26771_ (.A0(_07528_),
    .A1(_07834_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net244));
 sky130_fd_sc_hd__inv_1 _26772_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .Y(_07835_));
 sky130_fd_sc_hd__mux2i_1 _26773_ (.A0(_07522_),
    .A1(_07835_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net245));
 sky130_fd_sc_hd__nand2_1 _26774_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .Y(_07836_));
 sky130_fd_sc_hd__o21ai_0 _26775_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07517_),
    .B1(_07836_),
    .Y(net246));
 sky130_fd_sc_hd__inv_1 _26776_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .Y(_07837_));
 sky130_fd_sc_hd__mux2i_1 _26777_ (.A0(_07707_),
    .A1(_07837_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(net247));
 sky130_fd_sc_hd__a21oi_1 _26778_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .A2(net3554),
    .B1(_07801_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_1 _26779_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .Y(_07839_));
 sky130_fd_sc_hd__o21ai_0 _26780_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07838_),
    .B1(_07839_),
    .Y(net248));
 sky130_fd_sc_hd__inv_1 _26781_ (.A(_07071_),
    .Y(net249));
 sky130_fd_sc_hd__nand2b_1 _26782_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .B(net128),
    .Y(_07840_));
 sky130_fd_sc_hd__a22o_1 _26783_ (.A1(net95),
    .A2(net249),
    .B1(_07840_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 sky130_fd_sc_hd__a31oi_1 _26784_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net95),
    .A3(net249),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_07841_));
 sky130_fd_sc_hd__a21oi_1 _26785_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .B1(_07841_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 sky130_fd_sc_hd__nor2_4 _26786_ (.A(net95),
    .B(_07544_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ));
 sky130_fd_sc_hd__nor2_1 _26787_ (.A(net95),
    .B(_07071_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 sky130_fd_sc_hd__a21oi_1 _26788_ (.A1(net3742),
    .A2(_06339_),
    .B1(net3448),
    .Y(_07842_));
 sky130_fd_sc_hd__o2111ai_1 _26789_ (.A1(_12171_),
    .A2(_06375_),
    .B1(\id_stage_i.controller_i.instr_valid_i ),
    .C1(_10795_),
    .D1(_10978_),
    .Y(_07843_));
 sky130_fd_sc_hd__nand2_1 _26790_ (.A(net3554),
    .B(net3443),
    .Y(_07844_));
 sky130_fd_sc_hd__o21ai_0 _26791_ (.A1(_07842_),
    .A2(_07843_),
    .B1(_07844_),
    .Y(\if_stage_i.instr_valid_id_d ));
 sky130_fd_sc_hd__dfrtp_4 _26792_ (.D(_00010_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 _26793_ (.D(_00011_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 _26794_ (.D(_00012_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 _26795_ (.D(_00013_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfstp_1 _26796_ (.D(_00014_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .SET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_core_clock (.A(clk_i),
    .X(delaynet_0_core_clock));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__buf_4 _26799_ (.A(net251),
    .X(alert_minor_o));
 sky130_fd_sc_hd__buf_4 _26800_ (.A(net252),
    .X(data_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _26801_ (.A(net253),
    .X(data_addr_o[1]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__buf_4 _26832_ (.A(net254),
    .X(instr_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _26833_ (.A(net255),
    .X(instr_addr_o[1]));
 sky130_fd_sc_hd__dfrtp_1 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .Q(core_busy_q),
    .RESET_B(net3956),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dlxtn_1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00008_),
    .Q(\core_clock_gate_i.en_latch ),
    .GATE_N(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_00015_),
    .Q(\cs_registers_i.mcountinhibit_q[0] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_00016_),
    .Q(\cs_registers_i.mcountinhibit_q[2] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_00017_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_00018_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_00019_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_00020_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_00021_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_00022_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_00023_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_00024_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_00025_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_00026_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_00027_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_00028_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_00029_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_00030_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_00031_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_00032_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_00033_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_00034_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_00035_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_00036_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_00037_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_00038_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_00039_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_00040_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_00041_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_00042_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_00043_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_00044_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_00045_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_00046_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_00047_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_00048_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_00049_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_00050_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_00051_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_00052_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_00053_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_00054_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_00055_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_00056_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_00057_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_00058_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_00059_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_00060_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_00061_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_00062_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_00063_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_00064_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_00065_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_00066_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_00067_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_00068_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_00069_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_00070_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_00071_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_00072_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_00073_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_00074_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_00075_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_00076_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_00077_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_00078_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_00079_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_00080_),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_00081_),
    .Q(\cs_registers_i.mhpmcounter[1856] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_00082_),
    .Q(\cs_registers_i.mhpmcounter[1866] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_00083_),
    .Q(\cs_registers_i.mhpmcounter[1867] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_00084_),
    .Q(\cs_registers_i.mhpmcounter[1868] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_00085_),
    .Q(\cs_registers_i.mhpmcounter[1869] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_00086_),
    .Q(\cs_registers_i.mhpmcounter[1870] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_00087_),
    .Q(\cs_registers_i.mhpmcounter[1871] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_00088_),
    .Q(\cs_registers_i.mhpmcounter[1872] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_00089_),
    .Q(\cs_registers_i.mhpmcounter[1873] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_00090_),
    .Q(\cs_registers_i.mhpmcounter[1874] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_00091_),
    .Q(\cs_registers_i.mhpmcounter[1875] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_00092_),
    .Q(\cs_registers_i.mhpmcounter[1857] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_00093_),
    .Q(\cs_registers_i.mhpmcounter[1876] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_00094_),
    .Q(\cs_registers_i.mhpmcounter[1877] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_00095_),
    .Q(\cs_registers_i.mhpmcounter[1878] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_00096_),
    .Q(\cs_registers_i.mhpmcounter[1879] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_00097_),
    .Q(\cs_registers_i.mhpmcounter[1880] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_00098_),
    .Q(\cs_registers_i.mhpmcounter[1881] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_00099_),
    .Q(\cs_registers_i.mhpmcounter[1882] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_00100_),
    .Q(\cs_registers_i.mhpmcounter[1883] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_00101_),
    .Q(\cs_registers_i.mhpmcounter[1884] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_00102_),
    .Q(\cs_registers_i.mhpmcounter[1885] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_00103_),
    .Q(\cs_registers_i.mhpmcounter[1858] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_00104_),
    .Q(\cs_registers_i.mhpmcounter[1886] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_00105_),
    .Q(\cs_registers_i.mhpmcounter[1887] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_00106_),
    .Q(\cs_registers_i.mhpmcounter[1888] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_00107_),
    .Q(\cs_registers_i.mhpmcounter[1889] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_00108_),
    .Q(\cs_registers_i.mhpmcounter[1890] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_00109_),
    .Q(\cs_registers_i.mhpmcounter[1891] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_00110_),
    .Q(\cs_registers_i.mhpmcounter[1892] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_00111_),
    .Q(\cs_registers_i.mhpmcounter[1893] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_00112_),
    .Q(\cs_registers_i.mhpmcounter[1894] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_00113_),
    .Q(\cs_registers_i.mhpmcounter[1895] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_00114_),
    .Q(\cs_registers_i.mhpmcounter[1859] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_00115_),
    .Q(\cs_registers_i.mhpmcounter[1896] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_00116_),
    .Q(\cs_registers_i.mhpmcounter[1897] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_00117_),
    .Q(\cs_registers_i.mhpmcounter[1898] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_00118_),
    .Q(\cs_registers_i.mhpmcounter[1899] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_00119_),
    .Q(\cs_registers_i.mhpmcounter[1900] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_00120_),
    .Q(\cs_registers_i.mhpmcounter[1901] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_00121_),
    .Q(\cs_registers_i.mhpmcounter[1902] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_00122_),
    .Q(\cs_registers_i.mhpmcounter[1903] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_00123_),
    .Q(\cs_registers_i.mhpmcounter[1904] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_00124_),
    .Q(\cs_registers_i.mhpmcounter[1905] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_00125_),
    .Q(\cs_registers_i.mhpmcounter[1860] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_00126_),
    .Q(\cs_registers_i.mhpmcounter[1906] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_00127_),
    .Q(\cs_registers_i.mhpmcounter[1907] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_00128_),
    .Q(\cs_registers_i.mhpmcounter[1908] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_00129_),
    .Q(\cs_registers_i.mhpmcounter[1909] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_00130_),
    .Q(\cs_registers_i.mhpmcounter[1910] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_00131_),
    .Q(\cs_registers_i.mhpmcounter[1911] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_00132_),
    .Q(\cs_registers_i.mhpmcounter[1912] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_00133_),
    .Q(\cs_registers_i.mhpmcounter[1913] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_00134_),
    .Q(\cs_registers_i.mhpmcounter[1914] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_00135_),
    .Q(\cs_registers_i.mhpmcounter[1915] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_00136_),
    .Q(\cs_registers_i.mhpmcounter[1861] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_00137_),
    .Q(\cs_registers_i.mhpmcounter[1916] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_00138_),
    .Q(\cs_registers_i.mhpmcounter[1917] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_00139_),
    .Q(\cs_registers_i.mhpmcounter[1918] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_00140_),
    .Q(\cs_registers_i.mhpmcounter[1919] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_00141_),
    .Q(\cs_registers_i.mhpmcounter[1862] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_00142_),
    .Q(\cs_registers_i.mhpmcounter[1863] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_00143_),
    .Q(\cs_registers_i.mhpmcounter[1864] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_00144_),
    .Q(\cs_registers_i.mhpmcounter[1865] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P_  (.D(_00145_),
    .Q(\cs_registers_i.priv_mode_id_o[0] ),
    .SET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P_  (.D(_00146_),
    .Q(\cs_registers_i.priv_mode_id_o[1] ),
    .SET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P_  (.D(_00147_),
    .Q(\cs_registers_i.dcsr_q[0] ),
    .SET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00148_),
    .Q(\cs_registers_i.dcsr_q[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00149_),
    .Q(\cs_registers_i.dcsr_q[12] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00150_),
    .Q(\cs_registers_i.dcsr_q[13] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00151_),
    .Q(\cs_registers_i.dcsr_q[15] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P_  (.D(_00152_),
    .Q(\cs_registers_i.dcsr_q[1] ),
    .SET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00153_),
    .Q(\cs_registers_i.dcsr_q[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00154_),
    .Q(\cs_registers_i.dcsr_q[6] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00155_),
    .Q(\cs_registers_i.dcsr_q[7] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00156_),
    .Q(\cs_registers_i.dcsr_q[8] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00157_),
    .Q(\cs_registers_i.csr_depc_o[10] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00158_),
    .Q(\cs_registers_i.csr_depc_o[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00159_),
    .Q(\cs_registers_i.csr_depc_o[12] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00160_),
    .Q(\cs_registers_i.csr_depc_o[13] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00161_),
    .Q(\cs_registers_i.csr_depc_o[14] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00162_),
    .Q(\cs_registers_i.csr_depc_o[15] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00163_),
    .Q(\cs_registers_i.csr_depc_o[16] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00164_),
    .Q(\cs_registers_i.csr_depc_o[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00165_),
    .Q(\cs_registers_i.csr_depc_o[18] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00166_),
    .Q(\cs_registers_i.csr_depc_o[19] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00167_),
    .Q(\cs_registers_i.csr_depc_o[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00168_),
    .Q(\cs_registers_i.csr_depc_o[20] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00169_),
    .Q(\cs_registers_i.csr_depc_o[21] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00170_),
    .Q(\cs_registers_i.csr_depc_o[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00171_),
    .Q(\cs_registers_i.csr_depc_o[23] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00172_),
    .Q(\cs_registers_i.csr_depc_o[24] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00173_),
    .Q(\cs_registers_i.csr_depc_o[25] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00174_),
    .Q(\cs_registers_i.csr_depc_o[26] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00175_),
    .Q(\cs_registers_i.csr_depc_o[27] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00176_),
    .Q(\cs_registers_i.csr_depc_o[28] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00177_),
    .Q(\cs_registers_i.csr_depc_o[29] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00178_),
    .Q(\cs_registers_i.csr_depc_o[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00179_),
    .Q(\cs_registers_i.csr_depc_o[30] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00180_),
    .Q(\cs_registers_i.csr_depc_o[31] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00181_),
    .Q(\cs_registers_i.csr_depc_o[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00182_),
    .Q(\cs_registers_i.csr_depc_o[4] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00183_),
    .Q(\cs_registers_i.csr_depc_o[5] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00184_),
    .Q(\cs_registers_i.csr_depc_o[6] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00185_),
    .Q(\cs_registers_i.csr_depc_o[7] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00186_),
    .Q(\cs_registers_i.csr_depc_o[8] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00187_),
    .Q(\cs_registers_i.csr_depc_o[9] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00188_),
    .Q(\cs_registers_i.dscratch0_q[0] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00189_),
    .Q(\cs_registers_i.dscratch0_q[10] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00190_),
    .Q(\cs_registers_i.dscratch0_q[11] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00191_),
    .Q(\cs_registers_i.dscratch0_q[12] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00192_),
    .Q(\cs_registers_i.dscratch0_q[13] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00193_),
    .Q(\cs_registers_i.dscratch0_q[14] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00194_),
    .Q(\cs_registers_i.dscratch0_q[15] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00195_),
    .Q(\cs_registers_i.dscratch0_q[16] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00196_),
    .Q(\cs_registers_i.dscratch0_q[17] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00197_),
    .Q(\cs_registers_i.dscratch0_q[18] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00198_),
    .Q(\cs_registers_i.dscratch0_q[19] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00199_),
    .Q(\cs_registers_i.dscratch0_q[1] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00200_),
    .Q(\cs_registers_i.dscratch0_q[20] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00201_),
    .Q(\cs_registers_i.dscratch0_q[21] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00202_),
    .Q(\cs_registers_i.dscratch0_q[22] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00203_),
    .Q(\cs_registers_i.dscratch0_q[23] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00204_),
    .Q(\cs_registers_i.dscratch0_q[24] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00205_),
    .Q(\cs_registers_i.dscratch0_q[25] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00206_),
    .Q(\cs_registers_i.dscratch0_q[26] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00207_),
    .Q(\cs_registers_i.dscratch0_q[27] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00208_),
    .Q(\cs_registers_i.dscratch0_q[28] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00209_),
    .Q(\cs_registers_i.dscratch0_q[29] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00210_),
    .Q(\cs_registers_i.dscratch0_q[2] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00211_),
    .Q(\cs_registers_i.dscratch0_q[30] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00212_),
    .Q(\cs_registers_i.dscratch0_q[31] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00213_),
    .Q(\cs_registers_i.dscratch0_q[3] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00214_),
    .Q(\cs_registers_i.dscratch0_q[4] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00215_),
    .Q(\cs_registers_i.dscratch0_q[5] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00216_),
    .Q(\cs_registers_i.dscratch0_q[6] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00217_),
    .Q(\cs_registers_i.dscratch0_q[7] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00218_),
    .Q(\cs_registers_i.dscratch0_q[8] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00219_),
    .Q(\cs_registers_i.dscratch0_q[9] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00220_),
    .Q(\cs_registers_i.dscratch1_q[0] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00221_),
    .Q(\cs_registers_i.dscratch1_q[10] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00222_),
    .Q(\cs_registers_i.dscratch1_q[11] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00223_),
    .Q(\cs_registers_i.dscratch1_q[12] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00224_),
    .Q(\cs_registers_i.dscratch1_q[13] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00225_),
    .Q(\cs_registers_i.dscratch1_q[14] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00226_),
    .Q(\cs_registers_i.dscratch1_q[15] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00227_),
    .Q(\cs_registers_i.dscratch1_q[16] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00228_),
    .Q(\cs_registers_i.dscratch1_q[17] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00229_),
    .Q(\cs_registers_i.dscratch1_q[18] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00230_),
    .Q(\cs_registers_i.dscratch1_q[19] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00231_),
    .Q(\cs_registers_i.dscratch1_q[1] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00232_),
    .Q(\cs_registers_i.dscratch1_q[20] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00233_),
    .Q(\cs_registers_i.dscratch1_q[21] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00234_),
    .Q(\cs_registers_i.dscratch1_q[22] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00235_),
    .Q(\cs_registers_i.dscratch1_q[23] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00236_),
    .Q(\cs_registers_i.dscratch1_q[24] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00237_),
    .Q(\cs_registers_i.dscratch1_q[25] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00238_),
    .Q(\cs_registers_i.dscratch1_q[26] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00239_),
    .Q(\cs_registers_i.dscratch1_q[27] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00240_),
    .Q(\cs_registers_i.dscratch1_q[28] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00241_),
    .Q(\cs_registers_i.dscratch1_q[29] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00242_),
    .Q(\cs_registers_i.dscratch1_q[2] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00243_),
    .Q(\cs_registers_i.dscratch1_q[30] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00244_),
    .Q(\cs_registers_i.dscratch1_q[31] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00245_),
    .Q(\cs_registers_i.dscratch1_q[3] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00246_),
    .Q(\cs_registers_i.dscratch1_q[4] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00247_),
    .Q(\cs_registers_i.dscratch1_q[5] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00248_),
    .Q(\cs_registers_i.dscratch1_q[6] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00249_),
    .Q(\cs_registers_i.dscratch1_q[7] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00250_),
    .Q(\cs_registers_i.dscratch1_q[8] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00251_),
    .Q(\cs_registers_i.dscratch1_q[9] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00252_),
    .Q(\cs_registers_i.mcause_q[0] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00253_),
    .Q(\cs_registers_i.mcause_q[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00254_),
    .Q(\cs_registers_i.mcause_q[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00255_),
    .Q(\cs_registers_i.mcause_q[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00256_),
    .Q(\cs_registers_i.mcause_q[4] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00257_),
    .Q(\cs_registers_i.mcause_q[5] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00258_),
    .Q(\cs_registers_i.csr_mepc_o[0] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00259_),
    .Q(\cs_registers_i.csr_mepc_o[10] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00260_),
    .Q(\cs_registers_i.csr_mepc_o[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00261_),
    .Q(\cs_registers_i.csr_mepc_o[12] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00262_),
    .Q(\cs_registers_i.csr_mepc_o[13] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00263_),
    .Q(\cs_registers_i.csr_mepc_o[14] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00264_),
    .Q(\cs_registers_i.csr_mepc_o[15] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00265_),
    .Q(\cs_registers_i.csr_mepc_o[16] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00266_),
    .Q(\cs_registers_i.csr_mepc_o[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00267_),
    .Q(\cs_registers_i.csr_mepc_o[18] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00268_),
    .Q(\cs_registers_i.csr_mepc_o[19] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00269_),
    .Q(\cs_registers_i.csr_mepc_o[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00270_),
    .Q(\cs_registers_i.csr_mepc_o[20] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00271_),
    .Q(\cs_registers_i.csr_mepc_o[21] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00272_),
    .Q(\cs_registers_i.csr_mepc_o[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00273_),
    .Q(\cs_registers_i.csr_mepc_o[23] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00274_),
    .Q(\cs_registers_i.csr_mepc_o[24] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00275_),
    .Q(\cs_registers_i.csr_mepc_o[25] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00276_),
    .Q(\cs_registers_i.csr_mepc_o[26] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00277_),
    .Q(\cs_registers_i.csr_mepc_o[27] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00278_),
    .Q(\cs_registers_i.csr_mepc_o[28] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00279_),
    .Q(\cs_registers_i.csr_mepc_o[29] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00280_),
    .Q(\cs_registers_i.csr_mepc_o[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00281_),
    .Q(\cs_registers_i.csr_mepc_o[30] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00282_),
    .Q(\cs_registers_i.csr_mepc_o[31] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00283_),
    .Q(\cs_registers_i.csr_mepc_o[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00284_),
    .Q(\cs_registers_i.csr_mepc_o[4] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00285_),
    .Q(\cs_registers_i.csr_mepc_o[5] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00286_),
    .Q(\cs_registers_i.csr_mepc_o[6] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00287_),
    .Q(\cs_registers_i.csr_mepc_o[7] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00288_),
    .Q(\cs_registers_i.csr_mepc_o[8] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00289_),
    .Q(\cs_registers_i.csr_mepc_o[9] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00290_),
    .Q(\cs_registers_i.mie_q[0] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00291_),
    .Q(\cs_registers_i.mie_q[10] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00292_),
    .Q(\cs_registers_i.mie_q[11] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00293_),
    .Q(\cs_registers_i.mie_q[12] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00294_),
    .Q(\cs_registers_i.mie_q[13] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00295_),
    .Q(\cs_registers_i.mie_q[14] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00296_),
    .Q(\cs_registers_i.mie_q[15] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00297_),
    .Q(\cs_registers_i.mie_q[16] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00298_),
    .Q(\cs_registers_i.mie_q[17] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00299_),
    .Q(\cs_registers_i.mie_q[1] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00300_),
    .Q(\cs_registers_i.mie_q[2] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00301_),
    .Q(\cs_registers_i.mie_q[3] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00302_),
    .Q(\cs_registers_i.mie_q[4] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00303_),
    .Q(\cs_registers_i.mie_q[5] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00304_),
    .Q(\cs_registers_i.mie_q[6] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00305_),
    .Q(\cs_registers_i.mie_q[7] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00306_),
    .Q(\cs_registers_i.mie_q[8] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00307_),
    .Q(\cs_registers_i.mie_q[9] ),
    .RESET_B(net3979),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00308_),
    .Q(\cs_registers_i.mscratch_q[0] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00309_),
    .Q(\cs_registers_i.mscratch_q[10] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00310_),
    .Q(\cs_registers_i.mscratch_q[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00311_),
    .Q(\cs_registers_i.mscratch_q[12] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00312_),
    .Q(\cs_registers_i.mscratch_q[13] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00313_),
    .Q(\cs_registers_i.mscratch_q[14] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00314_),
    .Q(\cs_registers_i.mscratch_q[15] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00315_),
    .Q(\cs_registers_i.mscratch_q[16] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00316_),
    .Q(\cs_registers_i.mscratch_q[17] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00317_),
    .Q(\cs_registers_i.mscratch_q[18] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00318_),
    .Q(\cs_registers_i.mscratch_q[19] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00319_),
    .Q(\cs_registers_i.mscratch_q[1] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00320_),
    .Q(\cs_registers_i.mscratch_q[20] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00321_),
    .Q(\cs_registers_i.mscratch_q[21] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00322_),
    .Q(\cs_registers_i.mscratch_q[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00323_),
    .Q(\cs_registers_i.mscratch_q[23] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00324_),
    .Q(\cs_registers_i.mscratch_q[24] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00325_),
    .Q(\cs_registers_i.mscratch_q[25] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00326_),
    .Q(\cs_registers_i.mscratch_q[26] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00327_),
    .Q(\cs_registers_i.mscratch_q[27] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00328_),
    .Q(\cs_registers_i.mscratch_q[28] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00329_),
    .Q(\cs_registers_i.mscratch_q[29] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00330_),
    .Q(\cs_registers_i.mscratch_q[2] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00331_),
    .Q(\cs_registers_i.mscratch_q[30] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00332_),
    .Q(\cs_registers_i.mscratch_q[31] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00333_),
    .Q(\cs_registers_i.mscratch_q[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00334_),
    .Q(\cs_registers_i.mscratch_q[4] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00335_),
    .Q(\cs_registers_i.mscratch_q[5] ),
    .RESET_B(net3976),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00336_),
    .Q(\cs_registers_i.mscratch_q[6] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00337_),
    .Q(\cs_registers_i.mscratch_q[7] ),
    .RESET_B(net3974),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00338_),
    .Q(\cs_registers_i.mscratch_q[8] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00339_),
    .Q(\cs_registers_i.mscratch_q[9] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00340_),
    .Q(\cs_registers_i.mstack_cause_q[0] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00341_),
    .Q(\cs_registers_i.mstack_cause_q[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00342_),
    .Q(\cs_registers_i.mstack_cause_q[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00343_),
    .Q(\cs_registers_i.mstack_cause_q[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00344_),
    .Q(\cs_registers_i.mstack_cause_q[4] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00345_),
    .Q(\cs_registers_i.mstack_cause_q[5] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00346_),
    .Q(\cs_registers_i.mstack_q[0] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00347_),
    .Q(\cs_registers_i.mstack_q[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P_  (.D(_00348_),
    .Q(\cs_registers_i.mstack_q[2] ),
    .SET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00349_),
    .Q(\cs_registers_i.mstack_epc_q[0] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00350_),
    .Q(\cs_registers_i.mstack_epc_q[10] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00351_),
    .Q(\cs_registers_i.mstack_epc_q[11] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00352_),
    .Q(\cs_registers_i.mstack_epc_q[12] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00353_),
    .Q(\cs_registers_i.mstack_epc_q[13] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00354_),
    .Q(\cs_registers_i.mstack_epc_q[14] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00355_),
    .Q(\cs_registers_i.mstack_epc_q[15] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00356_),
    .Q(\cs_registers_i.mstack_epc_q[16] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00357_),
    .Q(\cs_registers_i.mstack_epc_q[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00358_),
    .Q(\cs_registers_i.mstack_epc_q[18] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00359_),
    .Q(\cs_registers_i.mstack_epc_q[19] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00360_),
    .Q(\cs_registers_i.mstack_epc_q[1] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00361_),
    .Q(\cs_registers_i.mstack_epc_q[20] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00362_),
    .Q(\cs_registers_i.mstack_epc_q[21] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00363_),
    .Q(\cs_registers_i.mstack_epc_q[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00364_),
    .Q(\cs_registers_i.mstack_epc_q[23] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00365_),
    .Q(\cs_registers_i.mstack_epc_q[24] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00366_),
    .Q(\cs_registers_i.mstack_epc_q[25] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00367_),
    .Q(\cs_registers_i.mstack_epc_q[26] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00368_),
    .Q(\cs_registers_i.mstack_epc_q[27] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00369_),
    .Q(\cs_registers_i.mstack_epc_q[28] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00370_),
    .Q(\cs_registers_i.mstack_epc_q[29] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00371_),
    .Q(\cs_registers_i.mstack_epc_q[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00372_),
    .Q(\cs_registers_i.mstack_epc_q[30] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00373_),
    .Q(\cs_registers_i.mstack_epc_q[31] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00374_),
    .Q(\cs_registers_i.mstack_epc_q[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00375_),
    .Q(\cs_registers_i.mstack_epc_q[4] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00376_),
    .Q(\cs_registers_i.mstack_epc_q[5] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00377_),
    .Q(\cs_registers_i.mstack_epc_q[6] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00378_),
    .Q(\cs_registers_i.mstack_epc_q[7] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00379_),
    .Q(\cs_registers_i.mstack_epc_q[8] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00380_),
    .Q(\cs_registers_i.mstack_epc_q[9] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00381_),
    .Q(\cs_registers_i.csr_mstatus_tw_o ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00382_),
    .Q(\cs_registers_i.mstatus_q[1] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0N_  (.D(_00383_),
    .Q(\cs_registers_i.mstatus_q[2] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0N_  (.D(_00384_),
    .Q(\cs_registers_i.mstatus_q[3] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1N_  (.D(_00385_),
    .Q(\cs_registers_i.mstatus_q[4] ),
    .SET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0N_  (.D(_00386_),
    .Q(\cs_registers_i.csr_mstatus_mie_o ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00387_),
    .Q(\cs_registers_i.mtval_q[0] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00388_),
    .Q(\cs_registers_i.mtval_q[10] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00389_),
    .Q(\cs_registers_i.mtval_q[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00390_),
    .Q(\cs_registers_i.mtval_q[12] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00391_),
    .Q(\cs_registers_i.mtval_q[13] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00392_),
    .Q(\cs_registers_i.mtval_q[14] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00393_),
    .Q(\cs_registers_i.mtval_q[15] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00394_),
    .Q(\cs_registers_i.mtval_q[16] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00395_),
    .Q(\cs_registers_i.mtval_q[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00396_),
    .Q(\cs_registers_i.mtval_q[18] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00397_),
    .Q(\cs_registers_i.mtval_q[19] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00398_),
    .Q(\cs_registers_i.mtval_q[1] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00399_),
    .Q(\cs_registers_i.mtval_q[20] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00400_),
    .Q(\cs_registers_i.mtval_q[21] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00401_),
    .Q(\cs_registers_i.mtval_q[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00402_),
    .Q(\cs_registers_i.mtval_q[23] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00403_),
    .Q(\cs_registers_i.mtval_q[24] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00404_),
    .Q(\cs_registers_i.mtval_q[25] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00405_),
    .Q(\cs_registers_i.mtval_q[26] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00406_),
    .Q(\cs_registers_i.mtval_q[27] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00407_),
    .Q(\cs_registers_i.mtval_q[28] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00408_),
    .Q(\cs_registers_i.mtval_q[29] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00409_),
    .Q(\cs_registers_i.mtval_q[2] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00410_),
    .Q(\cs_registers_i.mtval_q[30] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00411_),
    .Q(\cs_registers_i.mtval_q[31] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00412_),
    .Q(\cs_registers_i.mtval_q[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00413_),
    .Q(\cs_registers_i.mtval_q[4] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00414_),
    .Q(\cs_registers_i.mtval_q[5] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00415_),
    .Q(\cs_registers_i.mtval_q[6] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00416_),
    .Q(\cs_registers_i.mtval_q[7] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00417_),
    .Q(\cs_registers_i.mtval_q[8] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00418_),
    .Q(\cs_registers_i.mtval_q[9] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00419_),
    .Q(\cs_registers_i.csr_mtvec_o[10] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00420_),
    .Q(\cs_registers_i.csr_mtvec_o[11] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00421_),
    .Q(\cs_registers_i.csr_mtvec_o[12] ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00422_),
    .Q(\cs_registers_i.csr_mtvec_o[13] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00423_),
    .Q(\cs_registers_i.csr_mtvec_o[14] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00424_),
    .Q(\cs_registers_i.csr_mtvec_o[15] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00425_),
    .Q(\cs_registers_i.csr_mtvec_o[16] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00426_),
    .Q(\cs_registers_i.csr_mtvec_o[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00427_),
    .Q(\cs_registers_i.csr_mtvec_o[18] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00428_),
    .Q(\cs_registers_i.csr_mtvec_o[19] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00429_),
    .Q(\cs_registers_i.csr_mtvec_o[20] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00430_),
    .Q(\cs_registers_i.csr_mtvec_o[21] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00431_),
    .Q(\cs_registers_i.csr_mtvec_o[22] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00432_),
    .Q(\cs_registers_i.csr_mtvec_o[23] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00433_),
    .Q(\cs_registers_i.csr_mtvec_o[24] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00434_),
    .Q(\cs_registers_i.csr_mtvec_o[25] ),
    .RESET_B(net3973),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00435_),
    .Q(\cs_registers_i.csr_mtvec_o[26] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00436_),
    .Q(\cs_registers_i.csr_mtvec_o[27] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00437_),
    .Q(\cs_registers_i.csr_mtvec_o[28] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00438_),
    .Q(\cs_registers_i.csr_mtvec_o[29] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00439_),
    .Q(\cs_registers_i.csr_mtvec_o[30] ),
    .RESET_B(net3975),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00440_),
    .Q(\cs_registers_i.csr_mtvec_o[31] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00441_),
    .Q(\cs_registers_i.csr_mtvec_o[8] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00442_),
    .Q(\cs_registers_i.csr_mtvec_o[9] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_00443_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_00444_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_00445_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_00446_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_00447_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_00448_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfstp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .SET_B(net3953),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_00449_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_00450_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_00451_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_00452_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_00453_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_00454_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_00455_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_00456_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_00457_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_00458_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_00459_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_00460_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_00461_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_00462_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_00463_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_00464_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_00465_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_00466_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_00467_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_00468_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_00469_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_00470_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_00471_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_00472_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .RESET_B(net3977),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_00473_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_00474_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_00475_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_00476_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_00477_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_00478_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_00479_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_00480_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_00481_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_00482_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_00483_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_00484_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_00485_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_00486_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_00487_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_00488_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_00489_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_00490_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_00491_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_00492_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_00493_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_00494_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_00495_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_00496_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_00497_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_00498_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_00499_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_00500_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_00501_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_00502_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_00503_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_00504_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_00505_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_00506_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_00507_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_00508_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_00509_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_00510_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_00511_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_00512_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \fetch_enable_q$_DFFE_PN0P_  (.D(_00513_),
    .Q(fetch_enable_q),
    .RESET_B(net3956),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P_  (.D(_00514_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P_  (.D(_00515_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P_  (.D(_00516_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P_  (.D(_00517_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P_  (.D(_00518_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P_  (.D(_00519_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P_  (.D(_00520_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P_  (.D(_00521_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P_  (.D(_00522_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P_  (.D(_00523_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P_  (.D(_00524_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P_  (.D(_00525_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P_  (.D(_00526_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P_  (.D(_00527_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P_  (.D(_00528_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P_  (.D(_00529_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P_  (.D(_00530_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P_  (.D(_00531_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P_  (.D(_00532_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P_  (.D(_00533_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P_  (.D(_00534_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P_  (.D(_00535_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P_  (.D(_00536_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P_  (.D(_00537_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P_  (.D(_00538_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P_  (.D(_00539_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P_  (.D(_00540_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P_  (.D(_00541_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P_  (.D(_00542_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P_  (.D(_00543_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P_  (.D(_00544_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P_  (.D(_00545_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P_  (.D(_00546_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P_  (.D(_00547_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P_  (.D(_00548_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P_  (.D(_00549_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P_  (.D(_00550_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P_  (.D(_00551_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P_  (.D(_00552_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P_  (.D(_00553_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P_  (.D(_00554_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P_  (.D(_00555_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P_  (.D(_00556_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P_  (.D(_00557_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P_  (.D(_00558_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P_  (.D(_00559_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P_  (.D(_00560_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P_  (.D(_00561_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P_  (.D(_00562_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P_  (.D(_00563_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P_  (.D(_00564_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P_  (.D(_00565_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P_  (.D(_00566_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P_  (.D(_00567_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P_  (.D(_00568_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P_  (.D(_00569_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P_  (.D(_00570_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P_  (.D(_00571_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P_  (.D(_00572_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P_  (.D(_00573_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P_  (.D(_00574_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P_  (.D(_00575_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P_  (.D(_00576_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P_  (.D(_00577_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P_  (.D(_00578_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P_  (.D(_00579_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P_  (.D(_00580_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P_  (.D(_00581_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P_  (.D(_00582_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P_  (.D(_00583_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P_  (.D(_00584_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P_  (.D(_00585_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P_  (.D(_00586_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P_  (.D(_00587_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P_  (.D(_00588_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P_  (.D(_00589_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P_  (.D(_00590_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P_  (.D(_00591_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P_  (.D(_00592_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P_  (.D(_00593_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P_  (.D(_00594_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P_  (.D(_00595_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P_  (.D(_00596_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P_  (.D(_00597_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P_  (.D(_00598_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P_  (.D(_00599_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P_  (.D(_00600_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P_  (.D(_00601_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P_  (.D(_00602_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P_  (.D(_00603_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P_  (.D(_00604_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P_  (.D(_00605_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P_  (.D(_00606_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P_  (.D(_00607_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P_  (.D(_00608_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P_  (.D(_00609_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P_  (.D(_00610_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P_  (.D(_00611_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P_  (.D(_00612_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P_  (.D(_00613_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P_  (.D(_00614_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P_  (.D(_00615_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P_  (.D(_00616_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P_  (.D(_00617_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P_  (.D(_00618_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P_  (.D(_00619_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P_  (.D(_00620_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P_  (.D(_00621_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P_  (.D(_00622_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P_  (.D(_00623_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P_  (.D(_00624_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P_  (.D(_00625_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P_  (.D(_00626_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P_  (.D(_00627_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P_  (.D(_00628_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P_  (.D(_00629_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P_  (.D(_00630_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P_  (.D(_00631_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P_  (.D(_00632_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P_  (.D(_00633_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P_  (.D(_00634_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P_  (.D(_00635_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P_  (.D(_00636_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P_  (.D(_00637_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P_  (.D(_00638_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P_  (.D(_00639_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P_  (.D(_00640_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P_  (.D(_00641_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P_  (.D(_00642_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P_  (.D(_00643_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P_  (.D(_00644_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P_  (.D(_00645_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P_  (.D(_00646_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P_  (.D(_00647_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P_  (.D(_00648_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P_  (.D(_00649_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P_  (.D(_00650_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P_  (.D(_00651_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P_  (.D(_00652_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P_  (.D(_00653_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P_  (.D(_00654_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P_  (.D(_00655_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P_  (.D(_00656_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P_  (.D(_00657_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P_  (.D(_00658_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P_  (.D(_00659_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P_  (.D(_00660_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P_  (.D(_00661_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P_  (.D(_00662_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P_  (.D(_00663_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P_  (.D(_00664_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P_  (.D(_00665_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P_  (.D(_00666_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P_  (.D(_00667_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P_  (.D(_00668_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P_  (.D(_00669_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P_  (.D(_00670_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P_  (.D(_00671_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P_  (.D(_00672_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P_  (.D(_00673_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P_  (.D(_00674_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P_  (.D(_00675_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P_  (.D(_00676_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P_  (.D(_00677_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P_  (.D(_00678_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P_  (.D(_00679_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P_  (.D(_00680_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P_  (.D(_00681_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P_  (.D(_00682_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P_  (.D(_00683_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P_  (.D(_00684_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P_  (.D(_00685_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P_  (.D(_00686_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P_  (.D(_00687_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P_  (.D(_00688_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P_  (.D(_00689_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P_  (.D(_00690_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P_  (.D(_00691_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P_  (.D(_00692_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P_  (.D(_00693_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P_  (.D(_00694_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P_  (.D(_00695_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P_  (.D(_00696_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P_  (.D(_00697_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P_  (.D(_00698_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P_  (.D(_00699_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P_  (.D(_00700_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P_  (.D(_00701_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P_  (.D(_00702_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P_  (.D(_00703_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P_  (.D(_00704_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P_  (.D(_00705_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P_  (.D(_00706_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P_  (.D(_00707_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P_  (.D(_00708_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P_  (.D(_00709_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P_  (.D(_00710_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P_  (.D(_00711_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P_  (.D(_00712_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P_  (.D(_00713_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P_  (.D(_00714_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P_  (.D(_00715_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P_  (.D(_00716_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P_  (.D(_00717_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P_  (.D(_00718_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P_  (.D(_00719_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P_  (.D(_00720_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P_  (.D(_00721_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P_  (.D(_00722_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P_  (.D(_00723_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P_  (.D(_00724_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P_  (.D(_00725_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P_  (.D(_00726_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P_  (.D(_00727_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P_  (.D(_00728_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P_  (.D(_00729_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P_  (.D(_00730_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P_  (.D(_00731_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P_  (.D(_00732_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P_  (.D(_00733_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P_  (.D(_00734_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P_  (.D(_00735_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P_  (.D(_00736_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P_  (.D(_00737_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P_  (.D(_00738_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P_  (.D(_00739_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P_  (.D(_00740_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P_  (.D(_00741_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P_  (.D(_00742_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P_  (.D(_00743_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P_  (.D(_00744_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P_  (.D(_00745_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P_  (.D(_00746_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P_  (.D(_00747_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P_  (.D(_00748_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P_  (.D(_00749_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P_  (.D(_00750_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P_  (.D(_00751_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P_  (.D(_00752_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P_  (.D(_00753_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P_  (.D(_00754_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P_  (.D(_00755_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P_  (.D(_00756_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P_  (.D(_00757_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P_  (.D(_00758_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P_  (.D(_00759_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P_  (.D(_00760_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P_  (.D(_00761_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P_  (.D(_00762_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P_  (.D(_00763_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P_  (.D(_00764_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P_  (.D(_00765_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P_  (.D(_00766_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P_  (.D(_00767_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P_  (.D(_00768_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P_  (.D(_00769_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P_  (.D(_00770_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P_  (.D(_00771_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P_  (.D(_00772_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P_  (.D(_00773_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P_  (.D(_00774_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P_  (.D(_00775_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P_  (.D(_00776_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P_  (.D(_00777_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P_  (.D(_00778_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P_  (.D(_00779_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P_  (.D(_00780_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P_  (.D(_00781_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P_  (.D(_00782_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P_  (.D(_00783_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P_  (.D(_00784_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P_  (.D(_00785_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P_  (.D(_00786_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P_  (.D(_00787_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P_  (.D(_00788_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P_  (.D(_00789_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P_  (.D(_00790_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P_  (.D(_00791_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P_  (.D(_00792_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P_  (.D(_00793_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P_  (.D(_00794_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P_  (.D(_00795_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P_  (.D(_00796_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P_  (.D(_00797_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P_  (.D(_00798_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P_  (.D(_00799_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P_  (.D(_00800_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P_  (.D(_00801_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P_  (.D(_00802_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P_  (.D(_00803_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P_  (.D(_00804_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P_  (.D(_00805_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P_  (.D(_00806_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P_  (.D(_00807_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P_  (.D(_00808_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P_  (.D(_00809_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P_  (.D(_00810_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P_  (.D(_00811_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P_  (.D(_00812_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P_  (.D(_00813_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P_  (.D(_00814_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P_  (.D(_00815_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P_  (.D(_00816_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P_  (.D(_00817_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P_  (.D(_00818_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P_  (.D(_00819_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P_  (.D(_00820_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P_  (.D(_00821_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P_  (.D(_00822_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P_  (.D(_00823_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P_  (.D(_00824_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P_  (.D(_00825_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P_  (.D(_00826_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P_  (.D(_00827_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P_  (.D(_00828_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P_  (.D(_00829_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P_  (.D(_00830_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P_  (.D(_00831_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P_  (.D(_00832_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P_  (.D(_00833_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P_  (.D(_00834_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P_  (.D(_00835_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P_  (.D(_00836_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P_  (.D(_00837_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P_  (.D(_00838_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P_  (.D(_00839_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P_  (.D(_00840_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P_  (.D(_00841_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P_  (.D(_00842_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P_  (.D(_00843_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P_  (.D(_00844_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P_  (.D(_00845_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P_  (.D(_00846_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P_  (.D(_00847_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P_  (.D(_00848_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P_  (.D(_00849_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P_  (.D(_00850_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P_  (.D(_00851_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P_  (.D(_00852_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P_  (.D(_00853_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P_  (.D(_00854_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P_  (.D(_00855_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P_  (.D(_00856_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P_  (.D(_00857_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P_  (.D(_00858_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P_  (.D(_00859_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P_  (.D(_00860_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P_  (.D(_00861_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P_  (.D(_00862_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P_  (.D(_00863_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P_  (.D(_00864_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P_  (.D(_00865_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P_  (.D(_00866_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P_  (.D(_00867_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P_  (.D(_00868_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P_  (.D(_00869_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P_  (.D(_00870_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P_  (.D(_00871_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P_  (.D(_00872_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P_  (.D(_00873_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P_  (.D(_00874_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P_  (.D(_00875_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P_  (.D(_00876_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P_  (.D(_00877_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P_  (.D(_00878_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P_  (.D(_00879_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P_  (.D(_00880_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P_  (.D(_00881_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P_  (.D(_00882_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P_  (.D(_00883_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P_  (.D(_00884_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P_  (.D(_00885_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P_  (.D(_00886_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P_  (.D(_00887_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P_  (.D(_00888_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P_  (.D(_00889_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P_  (.D(_00890_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P_  (.D(_00891_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P_  (.D(_00892_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P_  (.D(_00893_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P_  (.D(_00894_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P_  (.D(_00895_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P_  (.D(_00896_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P_  (.D(_00897_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P_  (.D(_00898_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P_  (.D(_00899_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P_  (.D(_00900_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P_  (.D(_00901_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P_  (.D(_00902_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P_  (.D(_00903_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P_  (.D(_00904_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P_  (.D(_00905_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P_  (.D(_00906_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P_  (.D(_00907_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P_  (.D(_00908_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P_  (.D(_00909_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P_  (.D(_00910_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P_  (.D(_00911_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P_  (.D(_00912_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P_  (.D(_00913_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P_  (.D(_00914_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P_  (.D(_00915_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P_  (.D(_00916_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P_  (.D(_00917_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P_  (.D(_00918_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P_  (.D(_00919_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P_  (.D(_00920_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P_  (.D(_00921_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P_  (.D(_00922_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P_  (.D(_00923_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P_  (.D(_00924_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P_  (.D(_00925_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P_  (.D(_00926_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P_  (.D(_00927_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P_  (.D(_00928_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P_  (.D(_00929_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P_  (.D(_00930_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P_  (.D(_00931_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P_  (.D(_00932_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P_  (.D(_00933_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P_  (.D(_00934_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P_  (.D(_00935_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P_  (.D(_00936_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P_  (.D(_00937_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P_  (.D(_00938_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P_  (.D(_00939_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P_  (.D(_00940_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P_  (.D(_00941_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P_  (.D(_00942_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P_  (.D(_00943_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P_  (.D(_00944_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P_  (.D(_00945_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P_  (.D(_00946_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P_  (.D(_00947_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P_  (.D(_00948_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P_  (.D(_00949_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P_  (.D(_00950_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P_  (.D(_00951_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P_  (.D(_00952_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P_  (.D(_00953_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P_  (.D(_00954_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P_  (.D(_00955_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P_  (.D(_00956_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P_  (.D(_00957_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P_  (.D(_00958_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P_  (.D(_00959_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P_  (.D(_00960_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P_  (.D(_00961_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P_  (.D(_00962_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P_  (.D(_00963_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P_  (.D(_00964_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P_  (.D(_00965_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P_  (.D(_00966_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P_  (.D(_00967_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P_  (.D(_00968_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P_  (.D(_00969_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P_  (.D(_00970_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P_  (.D(_00971_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P_  (.D(_00972_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P_  (.D(_00973_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P_  (.D(_00974_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P_  (.D(_00975_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P_  (.D(_00976_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P_  (.D(_00977_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P_  (.D(_00978_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P_  (.D(_00979_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P_  (.D(_00980_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P_  (.D(_00981_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P_  (.D(_00982_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P_  (.D(_00983_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P_  (.D(_00984_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P_  (.D(_00985_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P_  (.D(_00986_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P_  (.D(_00987_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P_  (.D(_00988_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P_  (.D(_00989_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P_  (.D(_00990_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P_  (.D(_00991_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P_  (.D(_00992_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P_  (.D(_00993_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P_  (.D(_00994_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P_  (.D(_00995_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P_  (.D(_00996_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P_  (.D(_00997_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P_  (.D(_00998_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P_  (.D(_00999_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P_  (.D(_01000_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P_  (.D(_01001_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P_  (.D(_01002_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P_  (.D(_01003_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P_  (.D(_01004_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P_  (.D(_01005_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P_  (.D(_01006_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P_  (.D(_01007_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P_  (.D(_01008_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P_  (.D(_01009_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P_  (.D(_01010_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P_  (.D(_01011_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P_  (.D(_01012_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P_  (.D(_01013_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P_  (.D(_01014_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P_  (.D(_01015_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P_  (.D(_01016_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P_  (.D(_01017_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P_  (.D(_01018_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P_  (.D(_01019_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P_  (.D(_01020_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P_  (.D(_01021_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P_  (.D(_01022_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P_  (.D(_01023_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P_  (.D(_01024_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P_  (.D(_01025_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P_  (.D(_01026_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P_  (.D(_01027_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P_  (.D(_01028_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P_  (.D(_01029_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P_  (.D(_01030_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P_  (.D(_01031_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P_  (.D(_01032_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P_  (.D(_01033_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P_  (.D(_01034_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P_  (.D(_01035_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P_  (.D(_01036_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P_  (.D(_01037_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P_  (.D(_01038_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P_  (.D(_01039_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P_  (.D(_01040_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P_  (.D(_01041_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P_  (.D(_01042_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P_  (.D(_01043_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P_  (.D(_01044_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P_  (.D(_01045_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P_  (.D(_01046_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P_  (.D(_01047_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P_  (.D(_01048_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P_  (.D(_01049_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P_  (.D(_01050_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P_  (.D(_01051_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P_  (.D(_01052_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P_  (.D(_01053_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P_  (.D(_01054_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P_  (.D(_01055_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P_  (.D(_01056_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P_  (.D(_01057_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P_  (.D(_01058_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P_  (.D(_01059_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P_  (.D(_01060_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P_  (.D(_01061_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P_  (.D(_01062_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P_  (.D(_01063_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P_  (.D(_01064_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P_  (.D(_01065_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P_  (.D(_01066_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P_  (.D(_01067_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P_  (.D(_01068_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P_  (.D(_01069_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P_  (.D(_01070_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P_  (.D(_01071_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P_  (.D(_01072_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P_  (.D(_01073_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P_  (.D(_01074_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P_  (.D(_01075_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P_  (.D(_01076_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P_  (.D(_01077_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P_  (.D(_01078_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P_  (.D(_01079_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P_  (.D(_01080_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P_  (.D(_01081_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P_  (.D(_01082_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P_  (.D(_01083_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P_  (.D(_01084_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P_  (.D(_01085_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P_  (.D(_01086_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P_  (.D(_01087_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P_  (.D(_01088_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P_  (.D(_01089_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P_  (.D(_01090_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P_  (.D(_01091_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P_  (.D(_01092_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P_  (.D(_01093_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P_  (.D(_01094_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P_  (.D(_01095_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P_  (.D(_01096_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P_  (.D(_01097_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P_  (.D(_01098_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P_  (.D(_01099_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P_  (.D(_01100_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P_  (.D(_01101_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P_  (.D(_01102_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P_  (.D(_01103_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P_  (.D(_01104_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P_  (.D(_01105_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P_  (.D(_01106_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P_  (.D(_01107_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P_  (.D(_01108_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P_  (.D(_01109_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P_  (.D(_01110_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P_  (.D(_01111_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P_  (.D(_01112_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P_  (.D(_01113_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P_  (.D(_01114_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P_  (.D(_01115_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P_  (.D(_01116_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P_  (.D(_01117_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P_  (.D(_01118_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P_  (.D(_01119_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P_  (.D(_01120_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P_  (.D(_01121_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P_  (.D(_01122_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P_  (.D(_01123_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P_  (.D(_01124_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P_  (.D(_01125_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P_  (.D(_01126_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P_  (.D(_01127_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P_  (.D(_01128_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P_  (.D(_01129_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P_  (.D(_01130_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P_  (.D(_01131_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P_  (.D(_01132_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P_  (.D(_01133_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P_  (.D(_01134_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P_  (.D(_01135_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P_  (.D(_01136_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P_  (.D(_01137_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P_  (.D(_01138_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P_  (.D(_01139_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P_  (.D(_01140_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P_  (.D(_01141_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P_  (.D(_01142_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P_  (.D(_01143_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P_  (.D(_01144_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P_  (.D(_01145_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P_  (.D(_01146_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P_  (.D(_01147_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P_  (.D(_01148_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P_  (.D(_01149_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P_  (.D(_01150_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P_  (.D(_01151_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P_  (.D(_01152_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P_  (.D(_01153_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P_  (.D(_01154_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P_  (.D(_01155_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P_  (.D(_01156_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P_  (.D(_01157_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P_  (.D(_01158_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P_  (.D(_01159_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P_  (.D(_01160_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P_  (.D(_01161_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P_  (.D(_01162_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P_  (.D(_01163_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P_  (.D(_01164_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P_  (.D(_01165_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P_  (.D(_01166_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P_  (.D(_01167_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P_  (.D(_01168_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P_  (.D(_01169_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P_  (.D(_01170_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P_  (.D(_01171_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P_  (.D(_01172_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P_  (.D(_01173_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P_  (.D(_01174_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P_  (.D(_01175_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P_  (.D(_01176_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P_  (.D(_01177_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P_  (.D(_01178_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P_  (.D(_01179_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P_  (.D(_01180_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P_  (.D(_01181_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P_  (.D(_01182_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P_  (.D(_01183_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P_  (.D(_01184_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P_  (.D(_01185_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P_  (.D(_01186_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P_  (.D(_01187_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P_  (.D(_01188_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P_  (.D(_01189_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P_  (.D(_01190_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P_  (.D(_01191_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P_  (.D(_01192_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P_  (.D(_01193_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P_  (.D(_01194_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P_  (.D(_01195_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P_  (.D(_01196_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P_  (.D(_01197_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P_  (.D(_01198_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P_  (.D(_01199_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P_  (.D(_01200_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P_  (.D(_01201_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P_  (.D(_01202_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P_  (.D(_01203_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P_  (.D(_01204_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P_  (.D(_01205_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P_  (.D(_01206_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P_  (.D(_01207_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P_  (.D(_01208_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P_  (.D(_01209_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P_  (.D(_01210_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P_  (.D(_01211_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P_  (.D(_01212_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P_  (.D(_01213_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P_  (.D(_01214_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P_  (.D(_01215_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P_  (.D(_01216_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P_  (.D(_01217_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P_  (.D(_01218_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P_  (.D(_01219_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P_  (.D(_01220_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .RESET_B(net3970),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P_  (.D(_01221_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P_  (.D(_01222_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P_  (.D(_01223_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P_  (.D(_01224_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P_  (.D(_01225_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P_  (.D(_01226_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P_  (.D(_01227_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P_  (.D(_01228_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P_  (.D(_01229_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P_  (.D(_01230_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P_  (.D(_01231_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P_  (.D(_01232_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P_  (.D(_01233_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P_  (.D(_01234_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P_  (.D(_01235_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P_  (.D(_01236_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P_  (.D(_01237_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P_  (.D(_01238_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P_  (.D(_01239_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P_  (.D(_01240_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P_  (.D(_01241_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P_  (.D(_01242_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P_  (.D(_01243_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P_  (.D(_01244_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P_  (.D(_01245_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P_  (.D(_01246_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P_  (.D(_01247_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P_  (.D(_01248_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P_  (.D(_01249_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P_  (.D(_01250_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P_  (.D(_01251_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P_  (.D(_01252_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P_  (.D(_01253_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P_  (.D(_01254_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P_  (.D(_01255_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P_  (.D(_01256_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P_  (.D(_01257_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P_  (.D(_01258_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P_  (.D(_01259_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P_  (.D(_01260_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P_  (.D(_01261_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P_  (.D(_01262_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P_  (.D(_01263_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P_  (.D(_01264_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P_  (.D(_01265_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P_  (.D(_01266_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P_  (.D(_01267_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P_  (.D(_01268_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P_  (.D(_01269_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P_  (.D(_01270_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P_  (.D(_01271_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P_  (.D(_01272_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P_  (.D(_01273_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P_  (.D(_01274_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P_  (.D(_01275_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P_  (.D(_01276_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P_  (.D(_01277_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P_  (.D(_01278_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P_  (.D(_01279_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P_  (.D(_01280_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P_  (.D(_01281_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P_  (.D(_01282_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P_  (.D(_01283_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P_  (.D(_01284_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P_  (.D(_01285_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P_  (.D(_01286_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P_  (.D(_01287_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P_  (.D(_01288_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P_  (.D(_01289_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P_  (.D(_01290_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P_  (.D(_01291_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P_  (.D(_01292_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P_  (.D(_01293_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P_  (.D(_01294_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P_  (.D(_01295_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P_  (.D(_01296_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P_  (.D(_01297_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P_  (.D(_01298_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P_  (.D(_01299_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P_  (.D(_01300_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P_  (.D(_01301_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P_  (.D(_01302_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P_  (.D(_01303_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P_  (.D(_01304_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P_  (.D(_01305_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P_  (.D(_01306_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P_  (.D(_01307_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P_  (.D(_01308_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P_  (.D(_01309_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P_  (.D(_01310_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P_  (.D(_01311_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P_  (.D(_01312_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P_  (.D(_01313_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P_  (.D(_01314_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P_  (.D(_01315_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P_  (.D(_01316_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P_  (.D(_01317_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P_  (.D(_01318_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P_  (.D(_01319_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P_  (.D(_01320_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P_  (.D(_01321_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P_  (.D(_01322_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P_  (.D(_01323_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P_  (.D(_01324_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P_  (.D(_01325_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P_  (.D(_01326_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P_  (.D(_01327_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P_  (.D(_01328_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P_  (.D(_01329_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P_  (.D(_01330_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P_  (.D(_01331_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P_  (.D(_01332_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P_  (.D(_01333_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P_  (.D(_01334_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P_  (.D(_01335_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P_  (.D(_01336_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P_  (.D(_01337_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P_  (.D(_01338_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P_  (.D(_01339_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P_  (.D(_01340_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P_  (.D(_01341_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P_  (.D(_01342_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P_  (.D(_01343_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P_  (.D(_01344_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P_  (.D(_01345_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P_  (.D(_01346_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P_  (.D(_01347_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P_  (.D(_01348_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P_  (.D(_01349_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P_  (.D(_01350_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P_  (.D(_01351_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P_  (.D(_01352_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P_  (.D(_01353_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P_  (.D(_01354_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P_  (.D(_01355_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P_  (.D(_01356_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P_  (.D(_01357_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P_  (.D(_01358_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P_  (.D(_01359_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P_  (.D(_01360_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P_  (.D(_01361_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P_  (.D(_01362_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P_  (.D(_01363_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P_  (.D(_01364_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P_  (.D(_01365_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P_  (.D(_01366_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P_  (.D(_01367_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P_  (.D(_01368_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P_  (.D(_01369_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P_  (.D(_01370_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P_  (.D(_01371_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P_  (.D(_01372_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P_  (.D(_01373_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P_  (.D(_01374_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P_  (.D(_01375_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P_  (.D(_01376_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P_  (.D(_01377_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P_  (.D(_01378_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P_  (.D(_01379_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P_  (.D(_01380_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P_  (.D(_01381_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P_  (.D(_01382_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P_  (.D(_01383_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P_  (.D(_01384_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P_  (.D(_01385_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P_  (.D(_01386_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P_  (.D(_01387_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P_  (.D(_01388_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P_  (.D(_01389_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P_  (.D(_01390_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P_  (.D(_01391_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P_  (.D(_01392_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P_  (.D(_01393_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P_  (.D(_01394_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P_  (.D(_01395_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P_  (.D(_01396_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P_  (.D(_01397_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P_  (.D(_01398_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P_  (.D(_01399_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P_  (.D(_01400_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P_  (.D(_01401_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P_  (.D(_01402_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P_  (.D(_01403_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P_  (.D(_01404_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P_  (.D(_01405_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P_  (.D(_01406_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P_  (.D(_01407_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P_  (.D(_01408_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P_  (.D(_01409_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P_  (.D(_01410_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P_  (.D(_01411_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P_  (.D(_01412_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P_  (.D(_01413_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P_  (.D(_01414_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P_  (.D(_01415_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P_  (.D(_01416_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P_  (.D(_01417_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P_  (.D(_01418_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P_  (.D(_01419_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P_  (.D(_01420_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P_  (.D(_01421_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P_  (.D(_01422_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P_  (.D(_01423_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P_  (.D(_01424_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P_  (.D(_01425_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P_  (.D(_01426_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P_  (.D(_01427_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P_  (.D(_01428_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P_  (.D(_01429_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P_  (.D(_01430_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P_  (.D(_01431_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P_  (.D(_01432_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P_  (.D(_01433_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P_  (.D(_01434_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P_  (.D(_01435_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P_  (.D(_01436_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P_  (.D(_01437_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P_  (.D(_01438_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P_  (.D(_01439_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P_  (.D(_01440_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P_  (.D(_01441_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P_  (.D(_01442_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P_  (.D(_01443_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P_  (.D(_01444_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P_  (.D(_01445_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P_  (.D(_01446_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P_  (.D(_01447_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P_  (.D(_01448_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P_  (.D(_01449_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P_  (.D(_01450_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P_  (.D(_01451_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P_  (.D(_01452_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P_  (.D(_01453_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P_  (.D(_01454_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P_  (.D(_01455_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P_  (.D(_01456_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P_  (.D(_01457_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P_  (.D(_01458_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P_  (.D(_01459_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P_  (.D(_01460_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P_  (.D(_01461_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P_  (.D(_01462_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P_  (.D(_01463_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P_  (.D(_01464_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P_  (.D(_01465_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P_  (.D(_01466_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P_  (.D(_01467_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P_  (.D(_01468_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P_  (.D(_01469_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P_  (.D(_01470_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P_  (.D(_01471_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P_  (.D(_01472_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P_  (.D(_01473_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P_  (.D(_01474_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P_  (.D(_01475_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P_  (.D(_01476_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P_  (.D(_01477_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P_  (.D(_01478_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P_  (.D(_01479_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .RESET_B(net3964),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P_  (.D(_01480_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P_  (.D(_01481_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .RESET_B(net3966),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P_  (.D(_01482_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P_  (.D(_01483_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P_  (.D(_01484_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P_  (.D(_01485_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P_  (.D(_01486_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P_  (.D(_01487_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P_  (.D(_01488_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P_  (.D(_01489_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P_  (.D(_01490_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .RESET_B(net3965),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P_  (.D(_01491_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P_  (.D(_01492_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .RESET_B(net3958),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P_  (.D(_01493_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P_  (.D(_01494_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P_  (.D(_01495_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .RESET_B(net3959),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P_  (.D(_01496_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .RESET_B(net3960),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P_  (.D(_01497_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .RESET_B(net3962),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P_  (.D(_01498_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P_  (.D(_01499_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .RESET_B(net3967),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P_  (.D(_01500_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P_  (.D(_01501_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .RESET_B(net3969),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P_  (.D(_01502_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .RESET_B(net3963),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P_  (.D(_01503_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .RESET_B(net3957),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P_  (.D(_01504_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .RESET_B(net3961),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P_  (.D(_01505_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .RESET_B(net3968),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.branch_set$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .Q(\id_stage_i.branch_set ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_01506_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_01507_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_01508_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_01509_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P_  (.D(_01510_),
    .Q(\cs_registers_i.debug_mode_i ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .Q(\id_stage_i.controller_i.exc_req_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .Q(\id_stage_i.controller_i.illegal_insn_q ),
    .RESET_B(net3954),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_i ),
    .Q(\id_stage_i.controller_i.load_err_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P_  (.D(_01511_),
    .Q(\cs_registers_i.nmi_mode_i ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_i ),
    .Q(\id_stage_i.controller_i.store_err_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_01512_),
    .Q(\id_stage_i.id_fsm_q ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P_  (.D(_01513_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P_  (.D(_01514_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P_  (.D(_01515_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P_  (.D(_01516_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P_  (.D(_01517_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P_  (.D(_01518_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P_  (.D(_01519_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P_  (.D(_01520_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P_  (.D(_01521_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P_  (.D(_01522_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P_  (.D(_01523_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P_  (.D(_01524_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P_  (.D(_01525_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P_  (.D(_01526_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P_  (.D(_01527_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P_  (.D(_01528_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P_  (.D(_01529_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P_  (.D(_01530_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P_  (.D(_01531_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P_  (.D(_01532_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P_  (.D(_01533_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P_  (.D(_01534_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P_  (.D(_01535_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P_  (.D(_01536_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P_  (.D(_01537_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P_  (.D(_01538_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P_  (.D(_01539_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P_  (.D(_01540_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P_  (.D(_01541_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P_  (.D(_01542_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P_  (.D(_01543_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P_  (.D(_01544_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P_  (.D(_01545_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P_  (.D(_01546_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P_  (.D(_01547_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P_  (.D(_01548_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P_  (.D(_01549_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P_  (.D(_01550_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P_  (.D(_01551_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P_  (.D(_01552_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P_  (.D(_01553_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P_  (.D(_01554_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P_  (.D(_01555_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P_  (.D(_01556_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P_  (.D(_01557_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P_  (.D(_01558_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P_  (.D(_01559_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P_  (.D(_01560_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P_  (.D(_01561_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P_  (.D(_01562_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P_  (.D(_01563_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P_  (.D(_01564_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P_  (.D(_01565_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P_  (.D(_01566_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P_  (.D(_01567_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P_  (.D(_01568_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P_  (.D(_01569_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P_  (.D(_01570_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P_  (.D(_01571_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P_  (.D(_01572_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .RESET_B(net3978),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P_  (.D(_01573_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P_  (.D(_01574_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P_  (.D(_01575_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P_  (.D(_01576_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P_  (.D(_01577_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P_  (.D(_01578_),
    .Q(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .RESET_B(net3953),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .RESET_B(net148),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ),
    .DE(net3399),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(net94),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[0] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[11] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[12] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[13] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[16] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[18] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[19] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[20] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[2] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[21] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[22] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[23] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[24] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[25] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[26] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[29] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ),
    .DE(net3417),
    .Q(\cs_registers_i.pc_if_i[31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[4] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[6] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[8] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ),
    .DE(net3418),
    .Q(\cs_registers_i.pc_if_i[10] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ),
    .DE(net3399),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ),
    .DE(net3400),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ),
    .DE(net3400),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ),
    .DE(net3400),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ),
    .DE(net3400),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ),
    .DE(net3402),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ),
    .DE(net3400),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ),
    .DE(net3401),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(net96),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(net107),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(net118),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(net121),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(net122),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(net123),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(net124),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(net125),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(net126),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(net127),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(net97),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(net98),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(net99),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(net100),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(net101),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(net102),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(net103),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(net104),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(net105),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(net106),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(net108),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(net109),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(net110),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(net111),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(net112),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(net113),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(net114),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(net115),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(net116),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(net117),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(net119),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(net120),
    .DE(net3741),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(net219),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(net220),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(net221),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(net222),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(net223),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(net224),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(net225),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(net226),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(net227),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(net228),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(net229),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(net230),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(net231),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(net232),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(net233),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(net234),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(net235),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(net236),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(net237),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(net467),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(net239),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(net240),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(net241),
    .DE(net3517),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(net242),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(net243),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(net244),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(net245),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(net246),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(net247),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(net248),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .RESET_B(net148),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.illegal_instr_o ),
    .DE(net3441),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(\if_stage_i.fetch_err ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_01579_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.is_compressed_o ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(_10769_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[10] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_10862_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_10898_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_10867_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_10873_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_10879_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_10776_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[2] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[3] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(_10892_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[5] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[7] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_10850_),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[0]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[0] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[10]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[10] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[11]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[11] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[12]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[12] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[12] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[13]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[13] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[14]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[14] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[15]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[15] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[16]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[16] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[17]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[17] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[18]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[18] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[19]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[19] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[1]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[1] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[20]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[20] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[21]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[21] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[22]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[22] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[23]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[23] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[24]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[24] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[25]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[25] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[25] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[26]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[26] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[27]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[27] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[27] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[28]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[28] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[28] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[29]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[29] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[29] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[2]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[2] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[30]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[30] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[30] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[31]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[31] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[3]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[3] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[3] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[4]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[4] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[5]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[5] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[5] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[6]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[6] ),
    .DE(net3441),
    .Q(\id_stage_i.controller_i.instr_i[6] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[7]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[7] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[8]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[8] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_id_o[9]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[9] ),
    .DE(net3441),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.instr_valid_id_o$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .Q(\id_stage_i.controller_i.instr_valid_i ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[10] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[10] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[11] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[11] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[12] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[12] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[13] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[13] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[14] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[15] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[16] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[17] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[18] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[18] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[19] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[19] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(net3948),
    .DE(net3441),
    .Q(\cs_registers_i.pc_id_i[1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[20] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[20] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[21] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[21] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[22] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[22] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[23] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[24] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[24] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[25] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[25] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[26] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[26] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[27] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[28] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[29] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[29] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[2] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[2] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[30] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[31] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[31] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[3] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[4] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[5] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[6] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[6] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[7] ),
    .DE(net3443),
    .Q(\cs_registers_i.pc_id_i[7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[8] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[8] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[9] ),
    .DE(net3442),
    .Q(\cs_registers_i.pc_id_i[9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P_  (.D(_01580_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P_  (.D(_01581_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P_  (.D(_01582_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P_  (.D(_01583_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P_  (.D(_01584_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P_  (.D(_01585_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P_  (.D(_01586_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P_  (.D(_01587_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P_  (.D(_01588_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P_  (.D(_01589_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P_  (.D(_01590_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P_  (.D(_01591_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P_  (.D(_01592_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P_  (.D(_01593_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P_  (.D(_01594_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P_  (.D(_01595_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P_  (.D(_01596_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P_  (.D(_01597_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P_  (.D(_01598_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P_  (.D(_01599_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P_  (.D(_01600_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P_  (.D(_01601_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P_  (.D(_01602_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P_  (.D(_01603_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P_  (.D(_01604_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .RESET_B(net3952),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P_  (.D(_01605_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P_  (.D(_01606_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P_  (.D(_01607_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P_  (.D(_01608_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P_  (.D(_01609_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .RESET_B(net3951),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P_  (.D(_01610_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P_  (.D(_01611_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .RESET_B(net3955),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_01612_),
    .Q(\load_store_unit_i.data_sign_ext_q ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.data_type_q[1]$_DFF_PN0_  (.D(_00006_),
    .Q(\load_store_unit_i.data_type_q[1] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.data_type_q[2]$_DFF_PN0_  (.D(_00007_),
    .Q(\load_store_unit_i.data_type_q[2] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_01613_),
    .Q(\load_store_unit_i.data_we_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_01614_),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_01615_),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_01616_),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_01617_),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_01618_),
    .Q(\load_store_unit_i.lsu_err_q ),
    .RESET_B(net3956),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_01619_),
    .Q(\load_store_unit_i.rdata_offset_q[0] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_01620_),
    .Q(\load_store_unit_i.rdata_offset_q[1] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_01621_),
    .Q(\load_store_unit_i.rdata_q[0] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_01622_),
    .Q(\load_store_unit_i.rdata_q[10] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_01623_),
    .Q(\load_store_unit_i.rdata_q[11] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_01624_),
    .Q(\load_store_unit_i.rdata_q[12] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_01625_),
    .Q(\load_store_unit_i.rdata_q[13] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_01626_),
    .Q(\load_store_unit_i.rdata_q[14] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_01627_),
    .Q(\load_store_unit_i.rdata_q[15] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_01628_),
    .Q(\load_store_unit_i.rdata_q[16] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_01629_),
    .Q(\load_store_unit_i.rdata_q[17] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_01630_),
    .Q(\load_store_unit_i.rdata_q[18] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_01631_),
    .Q(\load_store_unit_i.rdata_q[19] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_01632_),
    .Q(\load_store_unit_i.rdata_q[1] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_01633_),
    .Q(\load_store_unit_i.rdata_q[20] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_01634_),
    .Q(\load_store_unit_i.rdata_q[21] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_01635_),
    .Q(\load_store_unit_i.rdata_q[22] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_01636_),
    .Q(\load_store_unit_i.rdata_q[23] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_01637_),
    .Q(\load_store_unit_i.rdata_q[2] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_01638_),
    .Q(\load_store_unit_i.rdata_q[3] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_01639_),
    .Q(\load_store_unit_i.rdata_q[4] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_01640_),
    .Q(\load_store_unit_i.rdata_q[5] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_01641_),
    .Q(\load_store_unit_i.rdata_q[6] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_01642_),
    .Q(\load_store_unit_i.rdata_q[7] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_01643_),
    .Q(\load_store_unit_i.rdata_q[8] ),
    .RESET_B(net3972),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_01644_),
    .Q(\load_store_unit_i.rdata_q[9] ),
    .RESET_B(net3971),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_3957 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(boot_addr_i[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(boot_addr_i[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(boot_addr_i[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(boot_addr_i[13]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(boot_addr_i[14]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(boot_addr_i[15]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(boot_addr_i[16]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(boot_addr_i[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(boot_addr_i[18]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(boot_addr_i[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(boot_addr_i[20]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(boot_addr_i[21]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(boot_addr_i[22]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(boot_addr_i[23]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(boot_addr_i[24]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(boot_addr_i[25]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(boot_addr_i[26]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(boot_addr_i[27]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(boot_addr_i[28]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(boot_addr_i[29]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(boot_addr_i[30]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(boot_addr_i[31]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(boot_addr_i[8]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(boot_addr_i[9]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(data_err_i),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(data_gnt_i),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(data_rdata_i[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(data_rdata_i[10]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(data_rdata_i[11]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(data_rdata_i[12]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(data_rdata_i[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(data_rdata_i[14]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(data_rdata_i[15]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(data_rdata_i[16]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(data_rdata_i[17]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(data_rdata_i[18]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(data_rdata_i[19]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(data_rdata_i[1]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(data_rdata_i[20]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(data_rdata_i[21]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(data_rdata_i[22]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(data_rdata_i[23]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(data_rdata_i[24]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(data_rdata_i[25]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(data_rdata_i[26]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(data_rdata_i[27]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(data_rdata_i[28]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(data_rdata_i[29]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(data_rdata_i[2]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(data_rdata_i[30]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(data_rdata_i[31]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(data_rdata_i[3]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(data_rdata_i[4]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(data_rdata_i[5]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(data_rdata_i[6]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(data_rdata_i[7]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(data_rdata_i[8]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(data_rdata_i[9]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(data_rvalid_i),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(debug_req_i),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(fetch_enable_i),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(hart_id_i[0]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(hart_id_i[10]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(hart_id_i[11]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(hart_id_i[12]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(hart_id_i[13]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(hart_id_i[14]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(hart_id_i[15]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(hart_id_i[16]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(hart_id_i[17]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(hart_id_i[18]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(hart_id_i[19]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(hart_id_i[1]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(hart_id_i[20]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(hart_id_i[21]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(hart_id_i[22]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(hart_id_i[23]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(hart_id_i[24]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(hart_id_i[25]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(hart_id_i[26]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(hart_id_i[27]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(hart_id_i[28]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(hart_id_i[29]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(hart_id_i[2]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(hart_id_i[30]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(hart_id_i[31]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(hart_id_i[3]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(hart_id_i[4]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(hart_id_i[5]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(hart_id_i[6]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(hart_id_i[7]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(hart_id_i[8]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(hart_id_i[9]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(instr_err_i),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(instr_gnt_i),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(instr_rdata_i[0]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(instr_rdata_i[10]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(instr_rdata_i[11]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(instr_rdata_i[12]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(instr_rdata_i[13]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(instr_rdata_i[14]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(instr_rdata_i[15]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(instr_rdata_i[16]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(instr_rdata_i[17]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(instr_rdata_i[18]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(instr_rdata_i[19]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(instr_rdata_i[1]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(instr_rdata_i[20]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(instr_rdata_i[21]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input110 (.A(instr_rdata_i[22]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(instr_rdata_i[23]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(instr_rdata_i[24]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(instr_rdata_i[25]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(instr_rdata_i[26]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(instr_rdata_i[27]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(instr_rdata_i[28]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(instr_rdata_i[29]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(instr_rdata_i[2]),
    .X(net118));
 sky130_fd_sc_hd__buf_1 input119 (.A(instr_rdata_i[30]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input120 (.A(instr_rdata_i[31]),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input121 (.A(instr_rdata_i[3]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input122 (.A(instr_rdata_i[4]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(instr_rdata_i[5]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(instr_rdata_i[6]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(instr_rdata_i[7]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(instr_rdata_i[8]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(instr_rdata_i[9]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(instr_rvalid_i),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input129 (.A(irq_external_i),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input130 (.A(irq_fast_i[0]),
    .X(net130));
 sky130_fd_sc_hd__buf_1 input131 (.A(irq_fast_i[10]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(irq_fast_i[11]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input133 (.A(irq_fast_i[12]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input134 (.A(irq_fast_i[13]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input135 (.A(irq_fast_i[14]),
    .X(net135));
 sky130_fd_sc_hd__buf_1 input136 (.A(irq_fast_i[1]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 input137 (.A(irq_fast_i[2]),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(irq_fast_i[3]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(irq_fast_i[4]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(irq_fast_i[5]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(irq_fast_i[6]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(irq_fast_i[7]),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(irq_fast_i[8]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(irq_fast_i[9]),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(irq_nm_i),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(irq_software_i),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(irq_timer_i),
    .X(net147));
 sky130_fd_sc_hd__buf_12 input148 (.A(rst_ni),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(test_en_i),
    .X(net149));
 sky130_fd_sc_hd__buf_1 output150 (.A(net150),
    .X(core_sleep_o));
 sky130_fd_sc_hd__buf_1 output151 (.A(net3515),
    .X(data_addr_o[10]));
 sky130_fd_sc_hd__buf_1 output152 (.A(net152),
    .X(data_addr_o[11]));
 sky130_fd_sc_hd__buf_1 output153 (.A(net3514),
    .X(data_addr_o[12]));
 sky130_fd_sc_hd__buf_1 output154 (.A(net154),
    .X(data_addr_o[13]));
 sky130_fd_sc_hd__buf_1 output155 (.A(net3513),
    .X(data_addr_o[14]));
 sky130_fd_sc_hd__buf_1 output156 (.A(net3507),
    .X(data_addr_o[15]));
 sky130_fd_sc_hd__buf_1 output157 (.A(net3506),
    .X(data_addr_o[16]));
 sky130_fd_sc_hd__buf_1 output158 (.A(net420),
    .X(data_addr_o[17]));
 sky130_fd_sc_hd__buf_1 output159 (.A(net159),
    .X(data_addr_o[18]));
 sky130_fd_sc_hd__buf_1 output160 (.A(net160),
    .X(data_addr_o[19]));
 sky130_fd_sc_hd__buf_1 output161 (.A(net452),
    .X(data_addr_o[20]));
 sky130_fd_sc_hd__buf_1 output162 (.A(net162),
    .X(data_addr_o[21]));
 sky130_fd_sc_hd__buf_1 output163 (.A(net3503),
    .X(data_addr_o[22]));
 sky130_fd_sc_hd__buf_1 output164 (.A(net164),
    .X(data_addr_o[23]));
 sky130_fd_sc_hd__buf_1 output165 (.A(net272),
    .X(data_addr_o[24]));
 sky130_fd_sc_hd__buf_1 output166 (.A(net3495),
    .X(data_addr_o[25]));
 sky130_fd_sc_hd__buf_1 output167 (.A(net167),
    .X(data_addr_o[26]));
 sky130_fd_sc_hd__buf_1 output168 (.A(net168),
    .X(data_addr_o[27]));
 sky130_fd_sc_hd__buf_1 output169 (.A(net169),
    .X(data_addr_o[28]));
 sky130_fd_sc_hd__buf_1 output170 (.A(net292),
    .X(data_addr_o[29]));
 sky130_fd_sc_hd__buf_1 output171 (.A(net3549),
    .X(data_addr_o[2]));
 sky130_fd_sc_hd__buf_1 output172 (.A(net3473),
    .X(data_addr_o[30]));
 sky130_fd_sc_hd__buf_1 output173 (.A(net173),
    .X(data_addr_o[31]));
 sky130_fd_sc_hd__buf_1 output174 (.A(net174),
    .X(data_addr_o[3]));
 sky130_fd_sc_hd__buf_1 output175 (.A(net3535),
    .X(data_addr_o[4]));
 sky130_fd_sc_hd__buf_1 output176 (.A(net3537),
    .X(data_addr_o[5]));
 sky130_fd_sc_hd__buf_1 output177 (.A(net177),
    .X(data_addr_o[6]));
 sky130_fd_sc_hd__buf_1 output178 (.A(net3530),
    .X(data_addr_o[7]));
 sky130_fd_sc_hd__buf_1 output179 (.A(net3519),
    .X(data_addr_o[8]));
 sky130_fd_sc_hd__buf_1 output180 (.A(net3520),
    .X(data_addr_o[9]));
 sky130_fd_sc_hd__buf_1 output181 (.A(net181),
    .X(data_be_o[0]));
 sky130_fd_sc_hd__buf_1 output182 (.A(net182),
    .X(data_be_o[1]));
 sky130_fd_sc_hd__buf_1 output183 (.A(net183),
    .X(data_be_o[2]));
 sky130_fd_sc_hd__buf_1 output184 (.A(net184),
    .X(data_be_o[3]));
 sky130_fd_sc_hd__buf_1 output185 (.A(net185),
    .X(data_req_o));
 sky130_fd_sc_hd__buf_1 output186 (.A(net186),
    .X(data_wdata_o[0]));
 sky130_fd_sc_hd__buf_1 output187 (.A(net187),
    .X(data_wdata_o[10]));
 sky130_fd_sc_hd__buf_1 output188 (.A(net188),
    .X(data_wdata_o[11]));
 sky130_fd_sc_hd__buf_1 output189 (.A(net189),
    .X(data_wdata_o[12]));
 sky130_fd_sc_hd__buf_1 output190 (.A(net190),
    .X(data_wdata_o[13]));
 sky130_fd_sc_hd__buf_1 output191 (.A(net191),
    .X(data_wdata_o[14]));
 sky130_fd_sc_hd__buf_1 output192 (.A(net192),
    .X(data_wdata_o[15]));
 sky130_fd_sc_hd__buf_1 output193 (.A(net193),
    .X(data_wdata_o[16]));
 sky130_fd_sc_hd__buf_1 output194 (.A(net194),
    .X(data_wdata_o[17]));
 sky130_fd_sc_hd__buf_1 output195 (.A(net195),
    .X(data_wdata_o[18]));
 sky130_fd_sc_hd__buf_1 output196 (.A(net196),
    .X(data_wdata_o[19]));
 sky130_fd_sc_hd__buf_1 output197 (.A(net197),
    .X(data_wdata_o[1]));
 sky130_fd_sc_hd__buf_1 output198 (.A(net198),
    .X(data_wdata_o[20]));
 sky130_fd_sc_hd__buf_1 output199 (.A(net199),
    .X(data_wdata_o[21]));
 sky130_fd_sc_hd__buf_1 output200 (.A(net200),
    .X(data_wdata_o[22]));
 sky130_fd_sc_hd__buf_1 output201 (.A(net201),
    .X(data_wdata_o[23]));
 sky130_fd_sc_hd__buf_1 output202 (.A(net202),
    .X(data_wdata_o[24]));
 sky130_fd_sc_hd__buf_1 output203 (.A(net203),
    .X(data_wdata_o[25]));
 sky130_fd_sc_hd__buf_1 output204 (.A(net204),
    .X(data_wdata_o[26]));
 sky130_fd_sc_hd__buf_1 output205 (.A(net205),
    .X(data_wdata_o[27]));
 sky130_fd_sc_hd__buf_1 output206 (.A(net206),
    .X(data_wdata_o[28]));
 sky130_fd_sc_hd__buf_1 output207 (.A(net207),
    .X(data_wdata_o[29]));
 sky130_fd_sc_hd__buf_1 output208 (.A(net208),
    .X(data_wdata_o[2]));
 sky130_fd_sc_hd__buf_1 output209 (.A(net209),
    .X(data_wdata_o[30]));
 sky130_fd_sc_hd__buf_1 output210 (.A(net210),
    .X(data_wdata_o[31]));
 sky130_fd_sc_hd__buf_1 output211 (.A(net211),
    .X(data_wdata_o[3]));
 sky130_fd_sc_hd__buf_1 output212 (.A(net212),
    .X(data_wdata_o[4]));
 sky130_fd_sc_hd__buf_1 output213 (.A(net213),
    .X(data_wdata_o[5]));
 sky130_fd_sc_hd__buf_1 output214 (.A(net214),
    .X(data_wdata_o[6]));
 sky130_fd_sc_hd__buf_1 output215 (.A(net215),
    .X(data_wdata_o[7]));
 sky130_fd_sc_hd__buf_1 output216 (.A(net216),
    .X(data_wdata_o[8]));
 sky130_fd_sc_hd__buf_1 output217 (.A(net217),
    .X(data_wdata_o[9]));
 sky130_fd_sc_hd__buf_1 output218 (.A(net218),
    .X(data_we_o));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(instr_addr_o[10]));
 sky130_fd_sc_hd__buf_1 output220 (.A(net220),
    .X(instr_addr_o[11]));
 sky130_fd_sc_hd__buf_1 output221 (.A(net221),
    .X(instr_addr_o[12]));
 sky130_fd_sc_hd__buf_1 output222 (.A(net222),
    .X(instr_addr_o[13]));
 sky130_fd_sc_hd__buf_1 output223 (.A(net223),
    .X(instr_addr_o[14]));
 sky130_fd_sc_hd__buf_1 output224 (.A(net224),
    .X(instr_addr_o[15]));
 sky130_fd_sc_hd__buf_4 output225 (.A(net225),
    .X(instr_addr_o[16]));
 sky130_fd_sc_hd__buf_1 output226 (.A(net226),
    .X(instr_addr_o[17]));
 sky130_fd_sc_hd__buf_4 output227 (.A(net227),
    .X(instr_addr_o[18]));
 sky130_fd_sc_hd__buf_1 output228 (.A(net228),
    .X(instr_addr_o[19]));
 sky130_fd_sc_hd__buf_1 output229 (.A(net229),
    .X(instr_addr_o[20]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(instr_addr_o[21]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(instr_addr_o[22]));
 sky130_fd_sc_hd__buf_1 output232 (.A(net232),
    .X(instr_addr_o[23]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(instr_addr_o[24]));
 sky130_fd_sc_hd__buf_1 output234 (.A(net234),
    .X(instr_addr_o[25]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(instr_addr_o[26]));
 sky130_fd_sc_hd__buf_1 output236 (.A(net236),
    .X(instr_addr_o[27]));
 sky130_fd_sc_hd__buf_1 output237 (.A(net237),
    .X(instr_addr_o[28]));
 sky130_fd_sc_hd__buf_6 output238 (.A(net238),
    .X(instr_addr_o[29]));
 sky130_fd_sc_hd__buf_1 output239 (.A(net239),
    .X(instr_addr_o[2]));
 sky130_fd_sc_hd__buf_6 output240 (.A(net240),
    .X(instr_addr_o[30]));
 sky130_fd_sc_hd__buf_6 output241 (.A(net241),
    .X(instr_addr_o[31]));
 sky130_fd_sc_hd__buf_1 output242 (.A(net242),
    .X(instr_addr_o[3]));
 sky130_fd_sc_hd__buf_1 output243 (.A(net243),
    .X(instr_addr_o[4]));
 sky130_fd_sc_hd__buf_1 output244 (.A(net244),
    .X(instr_addr_o[5]));
 sky130_fd_sc_hd__buf_1 output245 (.A(net245),
    .X(instr_addr_o[6]));
 sky130_fd_sc_hd__buf_1 output246 (.A(net246),
    .X(instr_addr_o[7]));
 sky130_fd_sc_hd__buf_1 output247 (.A(net247),
    .X(instr_addr_o[8]));
 sky130_fd_sc_hd__buf_1 output248 (.A(net248),
    .X(instr_addr_o[9]));
 sky130_fd_sc_hd__buf_1 output249 (.A(net249),
    .X(instr_req_o));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(data_rdata_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(data_rdata_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(boot_addr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(data_rdata_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(boot_addr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(boot_addr_i[17]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_1__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_1 rebuffer95 (.A(net349),
    .X(net350));
 sky130_fd_sc_hd__buf_1 rebuffer72 (.A(_08959_),
    .X(net327));
 sky130_fd_sc_hd__buf_1 rebuffer71 (.A(net325),
    .X(net326));
 sky130_fd_sc_hd__buf_1 rebuffer19 (.A(net273),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_2_core_clock (.A(delaynet_2_core_clock),
    .X(delaynet_3_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload48 (.A(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload47 (.A(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3496 (.A(_09812_),
    .X(net3496));
 sky130_fd_sc_hd__buf_12 place3630 (.A(_03122_),
    .X(net3630));
 sky130_fd_sc_hd__buf_1 place3617 (.A(_08890_),
    .X(net3617));
 sky130_fd_sc_hd__buf_1 place3633 (.A(_02655_),
    .X(net3633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3674 (.A(_10448_),
    .X(net3674));
 sky130_fd_sc_hd__buf_1 place3669 (.A(_03310_),
    .X(net3669));
 sky130_fd_sc_hd__buf_12 place3687 (.A(net373),
    .X(net3687));
 sky130_fd_sc_hd__buf_12 place3792 (.A(net413),
    .X(net3792));
 sky130_fd_sc_hd__buf_1 place3731 (.A(_03471_),
    .X(net3731));
 sky130_fd_sc_hd__buf_8 place3767 (.A(_08604_),
    .X(net3767));
 sky130_fd_sc_hd__buf_1 place3736 (.A(_08623_),
    .X(net3736));
 sky130_fd_sc_hd__buf_12 place3777 (.A(net258),
    .X(net3777));
 sky130_fd_sc_hd__buf_1 place3753 (.A(_07905_),
    .X(net3753));
 sky130_fd_sc_hd__buf_12 place3751 (.A(_07960_),
    .X(net3751));
 sky130_fd_sc_hd__buf_2 place3762 (.A(_08910_),
    .X(net3762));
 sky130_fd_sc_hd__buf_12 place3760 (.A(_01681_),
    .X(net3760));
 sky130_fd_sc_hd__clkbuf_2 place3766 (.A(net407),
    .X(net3766));
 sky130_fd_sc_hd__buf_12 place3764 (.A(_08829_),
    .X(net3764));
 sky130_fd_sc_hd__buf_12 place3773 (.A(net3772),
    .X(net3773));
 sky130_fd_sc_hd__buf_1 place3817 (.A(_07927_),
    .X(net3817));
 sky130_fd_sc_hd__buf_12 place3970 (.A(net3967),
    .X(net3970));
 sky130_fd_sc_hd__buf_6 place3900 (.A(net284),
    .X(net3900));
 sky130_fd_sc_hd__conb_1 _26832__5 (.LO(net254));
 sky130_fd_sc_hd__clkbuf_4 place3934 (.A(net3933),
    .X(net3934));
 sky130_fd_sc_hd__buf_16 place3873 (.A(net3859),
    .X(net3873));
 sky130_fd_sc_hd__buf_1 place3826 (.A(\cs_registers_i.pc_id_i[26] ),
    .X(net3826));
 sky130_fd_sc_hd__buf_12 place3912 (.A(net3908),
    .X(net3912));
 sky130_fd_sc_hd__buf_12 place3403 (.A(_04916_),
    .X(net3403));
 sky130_fd_sc_hd__conb_1 _26801__4 (.LO(net253));
 sky130_fd_sc_hd__buf_12 place3940 (.A(net356),
    .X(net3940));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_6__leaf_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload14 (.A(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload17 (.A(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload36 (.A(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload35 (.A(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3964 (.A(net3960),
    .X(net3964));
 sky130_fd_sc_hd__buf_12 place3937 (.A(net3936),
    .X(net3937));
 sky130_fd_sc_hd__buf_12 place3967 (.A(net148),
    .X(net3967));
 sky130_fd_sc_hd__buf_12 place3933 (.A(net396),
    .X(net3933));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__buf_6 place3932 (.A(net3931),
    .X(net3932));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__buf_4 place3907 (.A(net3906),
    .X(net3907));
 sky130_fd_sc_hd__buf_12 place3906 (.A(net318),
    .X(net3906));
 sky130_fd_sc_hd__buf_12 place3410 (.A(_04122_),
    .X(net3410));
 sky130_fd_sc_hd__clkinvlp_4 clkload34 (.A(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload33 (.A(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload32 (.A(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload31 (.A(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload24 (.A(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3922 (.A(net3917),
    .X(net3922));
 sky130_fd_sc_hd__buf_12 place3921 (.A(net346),
    .X(net3921));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3963 (.A(net3960),
    .X(net3963));
 sky130_fd_sc_hd__buf_12 place3969 (.A(net3968),
    .X(net3969));
 sky130_fd_sc_hd__buf_12 place3931 (.A(net396),
    .X(net3931));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__conb_1 _26799__2 (.LO(net251));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3966 (.A(net3960),
    .X(net3966));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3955 (.A(net3954),
    .X(net3955));
 sky130_fd_sc_hd__buf_12 place3872 (.A(net3867),
    .X(net3872));
 sky130_fd_sc_hd__buf_8 place3402 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .X(net3402));
 sky130_fd_sc_hd__buf_12 place3871 (.A(net3867),
    .X(net3871));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_0__leaf_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload30 (.A(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload21 (.A(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload23 (.A(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload20 (.A(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload29 (.A(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload28 (.A(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload22 (.A(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload27 (.A(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload25 (.A(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3949 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .X(net3949));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net3530));
 sky130_fd_sc_hd__buf_12 place3948 (.A(\cs_registers_i.pc_if_i[1] ),
    .X(net3948));
 sky130_fd_sc_hd__buf_1 place3643 (.A(_01775_),
    .X(net3643));
 sky130_fd_sc_hd__buf_1 place3950 (.A(\cs_registers_i.priv_mode_id_o[0] ),
    .X(net3950));
 sky130_fd_sc_hd__clkinv_8 clkload26 (.A(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3747 (.A(net3744),
    .X(net3747));
 sky130_fd_sc_hd__buf_12 place3441 (.A(net3440),
    .X(net3441));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_5__leaf_clk_i_regs));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_07617_));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_3_0__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_3_1__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3404 (.A(_04817_),
    .X(net3404));
 sky130_fd_sc_hd__buf_1 place3428 (.A(_11899_),
    .X(net3428));
 sky130_fd_sc_hd__clkinv_16 clkload5 (.A(clknet_3_6__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_4__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3405 (.A(_04701_),
    .X(net3405));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3426 (.A(_12049_),
    .X(net3426));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net3496));
 sky130_fd_sc_hd__buf_1 place3423 (.A(_04676_),
    .X(net3423));
 sky130_fd_sc_hd__buf_1 place3420 (.A(_07723_),
    .X(net3420));
 sky130_fd_sc_hd__buf_12 place3413 (.A(_03775_),
    .X(net3413));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_07683_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net3497));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net3497));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_08261_));
 sky130_fd_sc_hd__buf_12 place3951 (.A(net148),
    .X(net3951));
 sky130_fd_sc_hd__buf_12 place3947 (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(net3947));
 sky130_fd_sc_hd__buf_12 place3952 (.A(net3951),
    .X(net3952));
 sky130_fd_sc_hd__buf_12 place3953 (.A(net3952),
    .X(net3953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_3__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3746 (.A(net3745),
    .X(net3746));
 sky130_fd_sc_hd__buf_6 place3440 (.A(_00009_),
    .X(net3440));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(hart_id_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(data_rdata_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(data_rdata_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(data_rdata_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(data_rdata_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(data_rdata_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(data_rdata_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(hart_id_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(data_rdata_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\ex_block_i.alu_i.imd_val_q_i[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(hart_id_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(hart_id_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(hart_id_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net3693));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(rst_ni));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net3681));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(data_rdata_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(data_rdata_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(data_rdata_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(data_rdata_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_02679_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(data_rdata_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(data_rdata_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(data_rdata_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(data_rdata_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(data_rdata_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(data_rdata_i[20]));
 sky130_fd_sc_hd__buf_12 place3425 (.A(_03408_),
    .X(net3425));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload10 (.A(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3406 (.A(_04593_),
    .X(net3406));
 sky130_fd_sc_hd__buf_12 place3407 (.A(_04460_),
    .X(net3407));
 sky130_fd_sc_hd__buf_12 place3408 (.A(_04371_),
    .X(net3408));
 sky130_fd_sc_hd__buf_12 place3409 (.A(_04247_),
    .X(net3409));
 sky130_fd_sc_hd__buf_12 place3416 (.A(_03533_),
    .X(net3416));
 sky130_fd_sc_hd__buf_1 place3414 (.A(_07725_),
    .X(net3414));
 sky130_fd_sc_hd__buf_12 place3412 (.A(_03900_),
    .X(net3412));
 sky130_fd_sc_hd__buf_1 place3419 (.A(_07723_),
    .X(net3419));
 sky130_fd_sc_hd__buf_6 place3415 (.A(_04898_),
    .X(net3415));
 sky130_fd_sc_hd__buf_1 place3429 (.A(_04812_),
    .X(net3429));
 sky130_fd_sc_hd__buf_12 place3418 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .X(net3418));
 sky130_fd_sc_hd__buf_12 place3417 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .X(net3417));
 sky130_fd_sc_hd__buf_1 place3421 (.A(_07723_),
    .X(net3421));
 sky130_fd_sc_hd__buf_1 place3422 (.A(_04896_),
    .X(net3422));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(data_rdata_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(data_rdata_i[19]));
 sky130_fd_sc_hd__clkinv_4 clkload8 (.A(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3424 (.A(_04225_),
    .X(net3424));
 sky130_fd_sc_hd__buf_12 place3435 (.A(_11894_),
    .X(net3435));
 sky130_fd_sc_hd__buf_12 place3434 (.A(_11897_),
    .X(net3434));
 sky130_fd_sc_hd__clkinv_16 clkload6 (.A(clknet_3_7__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3427 (.A(_11924_),
    .X(net3427));
 sky130_fd_sc_hd__clkinv_16 clkload4 (.A(clknet_3_5__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload3 (.A(clknet_3_4__leaf_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_3__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3433 (.A(_03656_),
    .X(net3433));
 sky130_fd_sc_hd__buf_1 place3430 (.A(_04599_),
    .X(net3430));
 sky130_fd_sc_hd__buf_1 place3431 (.A(_04103_),
    .X(net3431));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(data_rdata_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(data_rdata_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(data_rdata_i[16]));
 sky130_fd_sc_hd__buf_12 place3442 (.A(net3440),
    .X(net3442));
 sky130_fd_sc_hd__buf_1 place3432 (.A(_03985_),
    .X(net3432));
 sky130_fd_sc_hd__buf_8 place3449 (.A(_10961_),
    .X(net3449));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_7__leaf_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3744 (.A(net321),
    .X(net3744));
 sky130_fd_sc_hd__buf_12 place3444 (.A(_04941_),
    .X(net3444));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_2__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .X(clknet_0_clk_i_regs));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(data_rdata_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(data_rdata_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(data_rdata_i[12]));
 sky130_fd_sc_hd__buf_12 place3447 (.A(_03090_),
    .X(net3447));
 sky130_fd_sc_hd__buf_1 place3445 (.A(_04596_),
    .X(net3445));
 sky130_fd_sc_hd__buf_1 place3448 (.A(_10961_),
    .X(net3448));
 sky130_fd_sc_hd__buf_12 place3741 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .X(net3741));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(boot_addr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(boot_addr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(boot_addr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net3519));
 sky130_fd_sc_hd__buf_12 place3446 (.A(_03232_),
    .X(net3446));
 sky130_fd_sc_hd__buf_12 place3745 (.A(net3744),
    .X(net3745));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_11270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_11270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net340));
 sky130_fd_sc_hd__clkbuf_2 place3723 (.A(net293),
    .X(net3723));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_09983_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_09721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_09583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net3530));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net3530));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net3486));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net3687));
 sky130_fd_sc_hd__buf_1 rebuffer220 (.A(_08307_),
    .X(net486));
 sky130_fd_sc_hd__buf_1 rebuffer219 (.A(_08307_),
    .X(net485));
 sky130_fd_sc_hd__buf_1 rebuffer218 (.A(_08669_),
    .X(net484));
 sky130_fd_sc_hd__buf_1 rebuffer217 (.A(_08619_),
    .X(net483));
 sky130_fd_sc_hd__buf_1 rebuffer215 (.A(net3473),
    .X(net481));
 sky130_fd_sc_hd__buf_1 rebuffer214 (.A(net3473),
    .X(net480));
 sky130_fd_sc_hd__buf_4 rebuffer213 (.A(_10489_),
    .X(net479));
 sky130_fd_sc_hd__buf_4 rebuffer208 (.A(_08884_),
    .X(net474));
 sky130_fd_sc_hd__buf_2 rebuffer207 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_1 rebuffer206 (.A(_08071_),
    .X(net472));
 sky130_fd_sc_hd__buf_1 rebuffer205 (.A(_08026_),
    .X(net471));
 sky130_fd_sc_hd__buf_1 rebuffer202 (.A(_10307_),
    .X(net468));
 sky130_fd_sc_hd__buf_1 rebuffer201 (.A(net238),
    .X(net467));
 sky130_fd_sc_hd__buf_1 rebuffer200 (.A(_07687_),
    .X(net466));
 sky130_fd_sc_hd__buf_1 rebuffer186 (.A(net161),
    .X(net452));
 sky130_fd_sc_hd__buf_1 rebuffer185 (.A(net161),
    .X(net451));
 sky130_fd_sc_hd__buf_1 rebuffer184 (.A(net447),
    .X(net450));
 sky130_fd_sc_hd__buf_1 rebuffer183 (.A(net447),
    .X(net449));
 sky130_fd_sc_hd__buf_1 rebuffer182 (.A(net447),
    .X(net448));
 sky130_fd_sc_hd__buf_6 rebuffer181 (.A(_01695_),
    .X(net447));
 sky130_fd_sc_hd__buf_8 rebuffer180 (.A(_01713_),
    .X(net446));
 sky130_fd_sc_hd__buf_1 rebuffer179 (.A(_01713_),
    .X(net445));
 sky130_fd_sc_hd__buf_1 rebuffer178 (.A(_01713_),
    .X(net444));
 sky130_fd_sc_hd__buf_6 rebuffer177 (.A(_01699_),
    .X(net443));
 sky130_fd_sc_hd__buf_1 rebuffer176 (.A(_01683_),
    .X(net442));
 sky130_fd_sc_hd__buf_1 rebuffer175 (.A(_07686_),
    .X(net441));
 sky130_fd_sc_hd__buf_1 rebuffer174 (.A(net3917),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_16 clone173 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_1 rebuffer172 (.A(net436),
    .X(net438));
 sky130_fd_sc_hd__buf_1 rebuffer171 (.A(net436),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__buf_8 rebuffer170 (.A(_09838_),
    .X(net436));
 sky130_fd_sc_hd__buf_1 rebuffer169 (.A(_08167_),
    .X(net435));
 sky130_fd_sc_hd__buf_12 rebuffer168 (.A(net3873),
    .X(net434));
 sky130_fd_sc_hd__buf_1 rebuffer167 (.A(_08578_),
    .X(net433));
 sky130_fd_sc_hd__buf_1 rebuffer166 (.A(net3712),
    .X(net432));
 sky130_fd_sc_hd__buf_2 rebuffer165 (.A(_08191_),
    .X(net431));
 sky130_fd_sc_hd__buf_2 rebuffer164 (.A(_07951_),
    .X(net430));
 sky130_fd_sc_hd__buf_1 rebuffer163 (.A(_07951_),
    .X(net429));
 sky130_fd_sc_hd__buf_1 rebuffer162 (.A(_07951_),
    .X(net428));
 sky130_fd_sc_hd__buf_1 rebuffer161 (.A(_07951_),
    .X(net427));
 sky130_fd_sc_hd__buf_1 rebuffer160 (.A(_07951_),
    .X(net426));
 sky130_fd_sc_hd__buf_1 rebuffer159 (.A(_08777_),
    .X(net425));
 sky130_fd_sc_hd__buf_1 rebuffer158 (.A(net3929),
    .X(net424));
 sky130_fd_sc_hd__buf_1 rebuffer157 (.A(net3929),
    .X(net423));
 sky130_fd_sc_hd__buf_1 rebuffer156 (.A(_09583_),
    .X(net422));
 sky130_fd_sc_hd__buf_1 rebuffer155 (.A(net158),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__buf_1 rebuffer153 (.A(_09536_),
    .X(net419));
 sky130_fd_sc_hd__buf_1 rebuffer152 (.A(_09785_),
    .X(net418));
 sky130_fd_sc_hd__mux2i_2 clone151 (.A0(net3707),
    .A1(net418),
    .S(_01681_),
    .Y(net417));
 sky130_fd_sc_hd__buf_1 rebuffer150 (.A(_08059_),
    .X(net416));
 sky130_fd_sc_hd__buf_2 rebuffer149 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_16 clone148 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__buf_4 rebuffer147 (.A(_08147_),
    .X(net413));
 sky130_fd_sc_hd__buf_12 place3459 (.A(_03278_),
    .X(net3459));
 sky130_fd_sc_hd__buf_2 rebuffer146 (.A(_08147_),
    .X(net412));
 sky130_fd_sc_hd__buf_1 rebuffer145 (.A(_08147_),
    .X(net411));
 sky130_fd_sc_hd__buf_2 rebuffer144 (.A(net409),
    .X(net410));
 sky130_fd_sc_hd__buf_6 rebuffer143 (.A(_09424_),
    .X(net409));
 sky130_fd_sc_hd__buf_1 rebuffer142 (.A(_08820_),
    .X(net408));
 sky130_fd_sc_hd__buf_6 rebuffer141 (.A(_08820_),
    .X(net407));
 sky130_fd_sc_hd__buf_1 rebuffer140 (.A(_09582_),
    .X(net406));
 sky130_fd_sc_hd__buf_1 rebuffer139 (.A(net414),
    .X(net405));
 sky130_fd_sc_hd__buf_2 rebuffer138 (.A(net3859),
    .X(net404));
 sky130_fd_sc_hd__buf_1 place3465 (.A(_03666_),
    .X(net3465));
 sky130_fd_sc_hd__buf_1 rebuffer137 (.A(net402),
    .X(net403));
 sky130_fd_sc_hd__buf_1 rebuffer136 (.A(_08798_),
    .X(net402));
 sky130_fd_sc_hd__buf_1 rebuffer135 (.A(_09211_),
    .X(net401));
 sky130_fd_sc_hd__buf_12 rebuffer134 (.A(_09093_),
    .X(net400));
 sky130_fd_sc_hd__buf_1 place3458 (.A(_04130_),
    .X(net3458));
 sky130_fd_sc_hd__buf_6 rebuffer133 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .X(net399));
 sky130_fd_sc_hd__buf_1 place3460 (.A(_02535_),
    .X(net3460));
 sky130_fd_sc_hd__buf_1 place3461 (.A(_10960_),
    .X(net3461));
 sky130_fd_sc_hd__buf_2 rebuffer132 (.A(_01680_),
    .X(net398));
 sky130_fd_sc_hd__buf_6 rebuffer131 (.A(_01680_),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_16 clone130 (.A(net399),
    .X(net396));
 sky130_fd_sc_hd__buf_6 rebuffer129 (.A(_07941_),
    .X(net395));
 sky130_fd_sc_hd__buf_1 rebuffer128 (.A(_08064_),
    .X(net394));
 sky130_fd_sc_hd__buf_1 place3462 (.A(_10957_),
    .X(net3462));
 sky130_fd_sc_hd__buf_1 rebuffer117 (.A(_08437_),
    .X(net393));
 sky130_fd_sc_hd__buf_1 rebuffer216 (.A(_08619_),
    .X(net482));
 sky130_fd_sc_hd__buf_6 rebuffer91 (.A(_07845_),
    .X(net391));
 sky130_fd_sc_hd__buf_1 rebuffer86 (.A(net389),
    .X(net390));
 sky130_fd_sc_hd__buf_12 rebuffer67 (.A(_09276_),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__buf_1 rebuffer54 (.A(_01710_),
    .X(net388));
 sky130_fd_sc_hd__buf_1 rebuffer48 (.A(_01710_),
    .X(net387));
 sky130_fd_sc_hd__buf_1 rebuffer40 (.A(net391),
    .X(net386));
 sky130_fd_sc_hd__buf_1 rebuffer39 (.A(_07845_),
    .X(net385));
 sky130_fd_sc_hd__o2111a_2 clone13 (.A1(_08003_),
    .A2(_08012_),
    .B1(_08049_),
    .C1(_08030_),
    .D1(_08037_),
    .X(net384));
 sky130_fd_sc_hd__buf_1 rebuffer12 (.A(_08050_),
    .X(net383));
 sky130_fd_sc_hd__buf_12 place3463 (.A(_05080_),
    .X(net3463));
 sky130_fd_sc_hd__buf_1 place3464 (.A(_04920_),
    .X(net3464));
 sky130_fd_sc_hd__buf_1 rebuffer7 (.A(_08094_),
    .X(net372));
 sky130_fd_sc_hd__buf_1 place3477 (.A(net3476),
    .X(net3477));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__buf_1 rebuffer127 (.A(_08436_),
    .X(net382));
 sky130_fd_sc_hd__buf_1 rebuffer126 (.A(_08057_),
    .X(net381));
 sky130_fd_sc_hd__buf_1 rebuffer125 (.A(_08057_),
    .X(net380));
 sky130_fd_sc_hd__buf_1 rebuffer124 (.A(\id_stage_i.controller_i.instr_i[25] ),
    .X(net379));
 sky130_fd_sc_hd__buf_6 rebuffer122 (.A(_07640_),
    .X(net377));
 sky130_fd_sc_hd__buf_1 rebuffer121 (.A(net375),
    .X(net376));
 sky130_fd_sc_hd__buf_6 rebuffer120 (.A(_08302_),
    .X(net375));
 sky130_fd_sc_hd__buf_1 place3466 (.A(_07580_),
    .X(net3466));
 sky130_fd_sc_hd__buf_6 rebuffer212 (.A(_08292_),
    .X(net478));
 sky130_fd_sc_hd__buf_6 rebuffer118 (.A(_09834_),
    .X(net373));
 sky130_fd_sc_hd__buf_1 rebuffer116 (.A(_08282_),
    .X(net371));
 sky130_fd_sc_hd__buf_6 rebuffer115 (.A(_08282_),
    .X(net370));
 sky130_fd_sc_hd__buf_6 rebuffer114 (.A(_09224_),
    .X(net369));
 sky130_fd_sc_hd__buf_1 rebuffer113 (.A(net367),
    .X(net368));
 sky130_fd_sc_hd__buf_1 place3468 (.A(_03421_),
    .X(net3468));
 sky130_fd_sc_hd__buf_6 rebuffer112 (.A(\id_stage_i.controller_i.instr_i[28] ),
    .X(net367));
 sky130_fd_sc_hd__buf_1 rebuffer111 (.A(\id_stage_i.controller_i.instr_i[28] ),
    .X(net366));
 sky130_fd_sc_hd__buf_12 place3471 (.A(net3470),
    .X(net3471));
 sky130_fd_sc_hd__buf_2 rebuffer110 (.A(_07945_),
    .X(net365));
 sky130_fd_sc_hd__buf_1 rebuffer109 (.A(_07945_),
    .X(net364));
 sky130_fd_sc_hd__buf_2 rebuffer108 (.A(_07945_),
    .X(net363));
 sky130_fd_sc_hd__buf_1 rebuffer107 (.A(_07945_),
    .X(net362));
 sky130_fd_sc_hd__buf_2 rebuffer106 (.A(_07945_),
    .X(net361));
 sky130_fd_sc_hd__buf_4 rebuffer105 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .X(net360));
 sky130_fd_sc_hd__bufbuf_16 clone104 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_6 rebuffer103 (.A(_07602_),
    .X(net358));
 sky130_fd_sc_hd__buf_1 rebuffer102 (.A(net356),
    .X(net357));
 sky130_fd_sc_hd__buf_8 rebuffer101 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net356));
 sky130_fd_sc_hd__buf_1 rebuffer100 (.A(\id_stage_i.controller_i.instr_i[30] ),
    .X(net355));
 sky130_fd_sc_hd__buf_1 rebuffer99 (.A(\id_stage_i.controller_i.instr_i[30] ),
    .X(net354));
 sky130_fd_sc_hd__buf_1 rebuffer98 (.A(_09219_),
    .X(net353));
 sky130_fd_sc_hd__buf_1 rebuffer97 (.A(net351),
    .X(net352));
 sky130_fd_sc_hd__buf_8 rebuffer96 (.A(_07987_),
    .X(net351));
 sky130_fd_sc_hd__buf_8 place3470 (.A(_10492_),
    .X(net3470));
 sky130_fd_sc_hd__buf_12 place3472 (.A(_02149_),
    .X(net3472));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__buf_6 rebuffer94 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .X(net349));
 sky130_fd_sc_hd__buf_4 rebuffer93 (.A(\id_stage_i.controller_i.instr_i[27] ),
    .X(net348));
 sky130_fd_sc_hd__buf_6 rebuffer92 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .X(net347));
 sky130_fd_sc_hd__bufbuf_16 clone91 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_8 rebuffer90 (.A(net395),
    .X(net345));
 sky130_fd_sc_hd__buf_2 rebuffer89 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net344));
 sky130_fd_sc_hd__buf_6 rebuffer88 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net343));
 sky130_fd_sc_hd__buf_12 rebuffer87 (.A(_08661_),
    .X(net342));
 sky130_fd_sc_hd__bufbuf_16 clone86 (.A(net344),
    .X(net341));
 sky130_fd_sc_hd__buf_8 rebuffer85 (.A(_08844_),
    .X(net340));
 sky130_fd_sc_hd__buf_1 rebuffer84 (.A(\id_stage_i.controller_i.instr_i[2] ),
    .X(net339));
 sky130_fd_sc_hd__buf_1 rebuffer83 (.A(\id_stage_i.controller_i.instr_i[2] ),
    .X(net338));
 sky130_fd_sc_hd__buf_1 rebuffer82 (.A(_07845_),
    .X(net337));
 sky130_fd_sc_hd__buf_1 rebuffer81 (.A(_08050_),
    .X(net336));
 sky130_fd_sc_hd__buf_1 rebuffer80 (.A(net384),
    .X(net335));
 sky130_fd_sc_hd__buf_2 rebuffer79 (.A(\id_stage_i.controller_i.instr_i[1] ),
    .X(net334));
 sky130_fd_sc_hd__buf_1 rebuffer78 (.A(_09062_),
    .X(net333));
 sky130_fd_sc_hd__buf_1 rebuffer77 (.A(net331),
    .X(net332));
 sky130_fd_sc_hd__buf_12 rebuffer76 (.A(_09452_),
    .X(net331));
 sky130_fd_sc_hd__buf_1 rebuffer75 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net330));
 sky130_fd_sc_hd__buf_6 rebuffer74 (.A(\id_stage_i.controller_i.instr_i[0] ),
    .X(net329));
 sky130_fd_sc_hd__buf_1 rebuffer73 (.A(_08959_),
    .X(net328));
 sky130_fd_sc_hd__buf_12 place3473 (.A(net172),
    .X(net3473));
 sky130_fd_sc_hd__buf_1 place3474 (.A(net170),
    .X(net3474));
 sky130_fd_sc_hd__clkbuf_2 place3476 (.A(_03115_),
    .X(net3476));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__buf_8 rebuffer70 (.A(\id_stage_i.controller_i.instr_i[4] ),
    .X(net325));
 sky130_fd_sc_hd__buf_1 rebuffer69 (.A(net343),
    .X(net324));
 sky130_fd_sc_hd__buf_1 rebuffer68 (.A(_10242_),
    .X(net323));
 sky130_fd_sc_hd__buf_1 place3478 (.A(_11685_),
    .X(net3478));
 sky130_fd_sc_hd__bufbuf_16 clone67 (.A(net324),
    .X(net322));
 sky130_fd_sc_hd__buf_6 rebuffer66 (.A(_08308_),
    .X(net321));
 sky130_fd_sc_hd__buf_1 rebuffer65 (.A(_08158_),
    .X(net320));
 sky130_fd_sc_hd__buf_1 rebuffer64 (.A(_08158_),
    .X(net319));
 sky130_fd_sc_hd__buf_1 rebuffer63 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net318));
 sky130_fd_sc_hd__buf_6 rebuffer62 (.A(_09153_),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 rebuffer61 (.A(_09151_),
    .X(net316));
 sky130_fd_sc_hd__buf_1 rebuffer60 (.A(_09151_),
    .X(net315));
 sky130_fd_sc_hd__buf_1 rebuffer59 (.A(_09151_),
    .X(net314));
 sky130_fd_sc_hd__buf_6 rebuffer58 (.A(_07976_),
    .X(net313));
 sky130_fd_sc_hd__buf_6 rebuffer57 (.A(_07976_),
    .X(net312));
 sky130_fd_sc_hd__buf_2 rebuffer56 (.A(_07976_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 rebuffer55 (.A(_09511_),
    .X(net310));
 sky130_fd_sc_hd__bufbuf_16 clone54 (.A(net346),
    .X(net309));
 sky130_fd_sc_hd__buf_1 rebuffer53 (.A(_08663_),
    .X(net308));
 sky130_fd_sc_hd__buf_6 rebuffer52 (.A(\id_stage_i.controller_i.instr_i[6] ),
    .X(net307));
 sky130_fd_sc_hd__buf_2 rebuffer51 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net306));
 sky130_fd_sc_hd__buf_1 rebuffer50 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net305));
 sky130_fd_sc_hd__buf_1 place3479 (.A(_11530_),
    .X(net3479));
 sky130_fd_sc_hd__buf_1 rebuffer49 (.A(_08754_),
    .X(net304));
 sky130_fd_sc_hd__bufbuf_16 clone48 (.A(net414),
    .X(net303));
 sky130_fd_sc_hd__buf_1 rebuffer47 (.A(_08488_),
    .X(net302));
 sky130_fd_sc_hd__buf_1 rebuffer46 (.A(_08660_),
    .X(net301));
 sky130_fd_sc_hd__buf_1 place3480 (.A(_11506_),
    .X(net3480));
 sky130_fd_sc_hd__buf_8 rebuffer45 (.A(_08095_),
    .X(net300));
 sky130_fd_sc_hd__buf_1 rebuffer44 (.A(_08095_),
    .X(net299));
 sky130_fd_sc_hd__buf_12 place3487 (.A(_10238_),
    .X(net3487));
 sky130_fd_sc_hd__buf_6 rebuffer43 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net298));
 sky130_fd_sc_hd__buf_2 rebuffer42 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net297));
 sky130_fd_sc_hd__buf_6 rebuffer41 (.A(_07941_),
    .X(net296));
 sky130_fd_sc_hd__buf_1 place3494 (.A(_11390_),
    .X(net3494));
 sky130_fd_sc_hd__buf_1 place3489 (.A(_02941_),
    .X(net3489));
 sky130_fd_sc_hd__bufbuf_16 clone40 (.A(net257),
    .X(net295));
 sky130_fd_sc_hd__bufbuf_16 clone39 (.A(net257),
    .X(net294));
 sky130_fd_sc_hd__buf_4 rebuffer38 (.A(_08197_),
    .X(net293));
 sky130_fd_sc_hd__buf_1 rebuffer37 (.A(net170),
    .X(net292));
 sky130_fd_sc_hd__buf_1 rebuffer36 (.A(_08242_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 rebuffer35 (.A(_08242_),
    .X(net290));
 sky130_fd_sc_hd__buf_1 rebuffer34 (.A(_08242_),
    .X(net289));
 sky130_fd_sc_hd__buf_1 rebuffer33 (.A(_08439_),
    .X(net288));
 sky130_fd_sc_hd__buf_6 rebuffer32 (.A(net286),
    .X(net287));
 sky130_fd_sc_hd__buf_6 rebuffer31 (.A(\id_stage_i.controller_i.instr_i[5] ),
    .X(net286));
 sky130_fd_sc_hd__buf_1 rebuffer30 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .X(net285));
 sky130_fd_sc_hd__buf_1 rebuffer29 (.A(net283),
    .X(net284));
 sky130_fd_sc_hd__buf_6 rebuffer28 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .X(net283));
 sky130_fd_sc_hd__buf_1 rebuffer27 (.A(_07999_),
    .X(net282));
 sky130_fd_sc_hd__buf_1 place3493 (.A(_11406_),
    .X(net3493));
 sky130_fd_sc_hd__buf_1 rebuffer25 (.A(net486),
    .X(net280));
 sky130_fd_sc_hd__buf_1 rebuffer24 (.A(net278),
    .X(net279));
 sky130_fd_sc_hd__buf_4 rebuffer23 (.A(_07987_),
    .X(net278));
 sky130_fd_sc_hd__buf_4 rebuffer22 (.A(_07987_),
    .X(net277));
 sky130_fd_sc_hd__buf_12 place3491 (.A(_11573_),
    .X(net3491));
 sky130_fd_sc_hd__clkbuf_2 rebuffer21 (.A(net351),
    .X(net276));
 sky130_fd_sc_hd__buf_1 rebuffer20 (.A(net351),
    .X(net275));
 sky130_fd_sc_hd__buf_1 place3492 (.A(_11426_),
    .X(net3492));
 sky130_fd_sc_hd__buf_12 place3514 (.A(net153),
    .X(net3514));
 sky130_fd_sc_hd__buf_12 place3498 (.A(_09252_),
    .X(net3498));
 sky130_fd_sc_hd__buf_12 place3500 (.A(_12010_),
    .X(net3500));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3499 (.A(_02640_),
    .X(net3499));
 sky130_fd_sc_hd__buf_12 rebuffer18 (.A(net165),
    .X(net273));
 sky130_fd_sc_hd__buf_1 rebuffer17 (.A(net165),
    .X(net272));
 sky130_fd_sc_hd__buf_6 rebuffer16 (.A(_07692_),
    .X(net271));
 sky130_fd_sc_hd__buf_1 rebuffer15 (.A(_08192_),
    .X(net270));
 sky130_fd_sc_hd__buf_2 rebuffer14 (.A(_08192_),
    .X(net269));
 sky130_fd_sc_hd__buf_1 rebuffer13 (.A(net342),
    .X(net268));
 sky130_fd_sc_hd__bufbuf_16 clone12 (.A(net346),
    .X(net267));
 sky130_fd_sc_hd__buf_6 rebuffer11 (.A(net263),
    .X(net266));
 sky130_fd_sc_hd__buf_1 rebuffer10 (.A(net263),
    .X(net265));
 sky130_fd_sc_hd__buf_2 rebuffer9 (.A(net263),
    .X(net264));
 sky130_fd_sc_hd__buf_12 rebuffer8 (.A(_08139_),
    .X(net263));
 sky130_fd_sc_hd__bufbuf_16 clone7 (.A(net359),
    .X(net262));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(_09019_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 rebuffer5 (.A(_08292_),
    .X(net260));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(_08292_),
    .X(net259));
 sky130_fd_sc_hd__buf_8 rebuffer3 (.A(net478),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__buf_6 rebuffer2 (.A(net256),
    .X(net257));
 sky130_fd_sc_hd__buf_8 rebuffer1 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_4_core_clock (.A(delaynet_4_core_clock),
    .X(clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_3_core_clock (.A(delaynet_3_core_clock),
    .X(delaynet_4_core_clock));
 sky130_fd_sc_hd__buf_2 place3502 (.A(_10027_),
    .X(net3502));
 sky130_fd_sc_hd__buf_12 place3504 (.A(_09945_),
    .X(net3504));
 sky130_fd_sc_hd__buf_1 place3505 (.A(net161),
    .X(net3505));
 sky130_fd_sc_hd__buf_12 place3506 (.A(net157),
    .X(net3506));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .X(delaynet_2_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .X(delaynet_1_core_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__inv_16 clkload176 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_8 clkload175 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload174 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_4 clkload173 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload172 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__inv_6 clkload171 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_8 clkload170 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__inv_6 clkload169 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_8 clkload168 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_8 clkload167 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinv_2 clkload166 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__bufinv_16 clkload165 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload164 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__buf_1 place3510 (.A(_02528_),
    .X(net3510));
 sky130_fd_sc_hd__inv_8 clkload163 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload162 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload161 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__inv_12 clkload160 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__buf_1 place3512 (.A(net421),
    .X(net3512));
 sky130_fd_sc_hd__clkinv_8 clkload159 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__buf_8 place3515 (.A(net151),
    .X(net3515));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload158 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinv_8 clkload157 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload156 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkinv_2 clkload155 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload154 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinv_8 clkload153 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__inv_12 clkload152 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__inv_8 clkload151 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_4 clkload150 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload149 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__inv_6 clkload148 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload147 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload146 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload145 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__buf_12 place3519 (.A(net179),
    .X(net3519));
 sky130_fd_sc_hd__clkinvlp_4 clkload144 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__bufinv_16 clkload143 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__inv_8 clkload142 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload141 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_2 clkload140 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_4 clkload139 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__buf_1 place3523 (.A(_01881_),
    .X(net3523));
 sky130_fd_sc_hd__bufinv_16 clkload138 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__inv_6 clkload137 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__buf_1 place3527 (.A(_11222_),
    .X(net3527));
 sky130_fd_sc_hd__inv_6 clkload136 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload135 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_4 clkload134 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__inv_4 clkload133 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_8 clkload132 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_8 clkload131 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__inv_12 clkload130 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__inv_8 clkload129 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__inv_6 clkload128 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__buf_1 place3521 (.A(_02283_),
    .X(net3521));
 sky130_fd_sc_hd__clkinvlp_4 clkload127 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload126 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__buf_1 place3526 (.A(_11661_),
    .X(net3526));
 sky130_fd_sc_hd__clkbuf_1 clkload125 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__inv_8 clkload124 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_4 clkload123 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload122 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload121 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__inv_12 clkload120 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__buf_12 place3524 (.A(_12755_),
    .X(net3524));
 sky130_fd_sc_hd__buf_1 place3525 (.A(_11723_),
    .X(net3525));
 sky130_fd_sc_hd__clkinv_8 clkload119 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__buf_1 place3528 (.A(_11142_),
    .X(net3528));
 sky130_fd_sc_hd__inv_6 clkload118 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3532 (.A(_12394_),
    .X(net3532));
 sky130_fd_sc_hd__inv_12 clkload117 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__buf_1 place3531 (.A(_01996_),
    .X(net3531));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__inv_12 clkload116 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_6 clkload115 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_8 clkload114 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__inv_12 clkload113 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__inv_12 clkload112 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload111 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_8 clkload110 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkinv_8 clkload109 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload108 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload107 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_8 clkload106 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_8 clkload105 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__inv_8 clkload104 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload103 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__inv_12 clkload101 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__inv_12 clkload100 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_2 clkload99 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_16 clkload98 (.A(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload97 (.A(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload96 (.A(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkinv_16 clkload95 (.A(clknet_3_4_0_clk));
 sky130_fd_sc_hd__inv_6 clkload94 (.A(clknet_3_3_0_clk));
 sky130_fd_sc_hd__inv_6 clkload93 (.A(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload92 (.A(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__buf_6 place3541 (.A(net304),
    .X(net3541));
 sky130_fd_sc_hd__buf_1 place3535 (.A(net175),
    .X(net3535));
 sky130_fd_sc_hd__buf_12 place3538 (.A(_10625_),
    .X(net3538));
 sky130_fd_sc_hd__buf_12 place3539 (.A(_10619_),
    .X(net3539));
 sky130_fd_sc_hd__buf_1 place3542 (.A(_02777_),
    .X(net3542));
 sky130_fd_sc_hd__buf_12 place3540 (.A(_10591_),
    .X(net3540));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3548 (.A(_11057_),
    .X(net3548));
 sky130_fd_sc_hd__buf_1 place3553 (.A(_08745_),
    .X(net3553));
 sky130_fd_sc_hd__buf_12 place3555 (.A(_06999_),
    .X(net3555));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__buf_12 place3554 (.A(_07494_),
    .X(net3554));
 sky130_fd_sc_hd__buf_12 place3556 (.A(_06418_),
    .X(net3556));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__buf_12 place3564 (.A(_12174_),
    .X(net3564));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__buf_12 place3558 (.A(_02051_),
    .X(net3558));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__buf_1 place3561 (.A(_01837_),
    .X(net3561));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__buf_12 place3562 (.A(_13118_),
    .X(net3562));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__buf_1 place3566 (.A(_11076_),
    .X(net3566));
 sky130_fd_sc_hd__buf_12 place3567 (.A(_10826_),
    .X(net3567));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3571 (.A(_03575_),
    .X(net3571));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__buf_1 place3569 (.A(_07520_),
    .X(net3569));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__buf_12 place3611 (.A(_12181_),
    .X(net3611));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_6 clkload91 (.A(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload90 (.A(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload89 (.A(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload88 (.A(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload87 (.A(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload86 (.A(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload85 (.A(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload84 (.A(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload83 (.A(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload82 (.A(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload81 (.A(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload80 (.A(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload79 (.A(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload78 (.A(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload77 (.A(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload76 (.A(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload75 (.A(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload74 (.A(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload73 (.A(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload72 (.A(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload71 (.A(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload70 (.A(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__clkinv_8 clkload69 (.A(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload68 (.A(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload67 (.A(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload65 (.A(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload64 (.A(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3575 (.A(_10701_),
    .X(net3575));
 sky130_fd_sc_hd__inv_6 clkload63 (.A(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload61 (.A(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload60 (.A(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload58 (.A(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload57 (.A(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload56 (.A(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload55 (.A(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload54 (.A(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload53 (.A(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload52 (.A(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload51 (.A(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload50 (.A(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3576 (.A(_08670_),
    .X(net3576));
 sky130_fd_sc_hd__inv_6 clkload49 (.A(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload46 (.A(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload45 (.A(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload44 (.A(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload43 (.A(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload42 (.A(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload41 (.A(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__clkinv_4 clkload40 (.A(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__buf_2 place3876 (.A(net3859),
    .X(net3876));
 sky130_fd_sc_hd__clkbuf_8 clkload39 (.A(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3580 (.A(_10610_),
    .X(net3580));
 sky130_fd_sc_hd__buf_1 place3877 (.A(net359),
    .X(net3877));
 sky130_fd_sc_hd__buf_6 place3879 (.A(net414),
    .X(net3879));
 sky130_fd_sc_hd__inv_8 clkload38 (.A(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__inv_8 clkload37 (.A(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3411 (.A(_03999_),
    .X(net3411));
 sky130_fd_sc_hd__buf_1 place3436 (.A(net3435),
    .X(net3436));
 sky130_fd_sc_hd__buf_12 place3870 (.A(net3867),
    .X(net3870));
 sky130_fd_sc_hd__buf_2 place3869 (.A(net3868),
    .X(net3869));
 sky130_fd_sc_hd__buf_8 place3437 (.A(net3435),
    .X(net3437));
 sky130_fd_sc_hd__buf_12 place3868 (.A(net3867),
    .X(net3868));
 sky130_fd_sc_hd__buf_12 place3438 (.A(net3435),
    .X(net3438));
 sky130_fd_sc_hd__buf_12 place3439 (.A(net3435),
    .X(net3439));
 sky130_fd_sc_hd__buf_12 place3878 (.A(net404),
    .X(net3878));
 sky130_fd_sc_hd__buf_1 place3857 (.A(net256),
    .X(net3857));
 sky130_fd_sc_hd__buf_12 place3401 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .X(net3401));
 sky130_fd_sc_hd__buf_1 place3399 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .X(net3399));
 sky130_fd_sc_hd__buf_6 place3400 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .X(net3400));
 sky130_fd_sc_hd__buf_12 place3914 (.A(net3913),
    .X(net3914));
 sky130_fd_sc_hd__buf_12 place3913 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net3913));
 sky130_fd_sc_hd__buf_12 place3896 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .X(net3896));
 sky130_fd_sc_hd__buf_12 place3978 (.A(net3977),
    .X(net3978));
 sky130_fd_sc_hd__buf_12 place3977 (.A(net3974),
    .X(net3977));
 sky130_fd_sc_hd__buf_16 place3884 (.A(net343),
    .X(net3884));
 sky130_fd_sc_hd__buf_4 place3883 (.A(net3882),
    .X(net3883));
 sky130_fd_sc_hd__buf_1 place3862 (.A(net3861),
    .X(net3862));
 sky130_fd_sc_hd__buf_12 place3850 (.A(net257),
    .X(net3850));
 sky130_fd_sc_hd__buf_12 place3851 (.A(net295),
    .X(net3851));
 sky130_fd_sc_hd__buf_6 place3853 (.A(net3852),
    .X(net3853));
 sky130_fd_sc_hd__buf_1 place3787 (.A(_08171_),
    .X(net3787));
 sky130_fd_sc_hd__buf_2 place3776 (.A(_08292_),
    .X(net3776));
 sky130_fd_sc_hd__buf_2 place3765 (.A(_08820_),
    .X(net3765));
 sky130_fd_sc_hd__buf_1 place3763 (.A(_08834_),
    .X(net3763));
 sky130_fd_sc_hd__buf_1 place3759 (.A(_01681_),
    .X(net3759));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3758 (.A(_01685_),
    .X(net3758));
 sky130_fd_sc_hd__buf_1 place3750 (.A(_08188_),
    .X(net3750));
 sky130_fd_sc_hd__buf_12 place3774 (.A(_08299_),
    .X(net3774));
 sky130_fd_sc_hd__buf_12 place3756 (.A(_07857_),
    .X(net3756));
 sky130_fd_sc_hd__buf_12 place3737 (.A(_08498_),
    .X(net3737));
 sky130_fd_sc_hd__buf_1 place3735 (.A(_09651_),
    .X(net3735));
 sky130_fd_sc_hd__buf_1 place3733 (.A(_10866_),
    .X(net3733));
 sky130_fd_sc_hd__buf_1 place3730 (.A(_06488_),
    .X(net3730));
 sky130_fd_sc_hd__buf_12 place3728 (.A(_07888_),
    .X(net3728));
 sky130_fd_sc_hd__buf_12 place3713 (.A(_08542_),
    .X(net3713));
 sky130_fd_sc_hd__buf_1 place3588 (.A(_09520_),
    .X(net3588));
 sky130_fd_sc_hd__buf_12 place3581 (.A(_10584_),
    .X(net3581));
 sky130_fd_sc_hd__buf_1 place3705 (.A(_08881_),
    .X(net3705));
 sky130_fd_sc_hd__buf_1 place3780 (.A(net371),
    .X(net3780));
 sky130_fd_sc_hd__buf_12 place3732 (.A(_03471_),
    .X(net3732));
 sky130_fd_sc_hd__buf_1 place3725 (.A(_08079_),
    .X(net3725));
 sky130_fd_sc_hd__buf_8 place3700 (.A(net314),
    .X(net3700));
 sky130_fd_sc_hd__buf_12 place3779 (.A(_08282_),
    .X(net3779));
 sky130_fd_sc_hd__buf_12 place3695 (.A(_09362_),
    .X(net3695));
 sky130_fd_sc_hd__buf_1 place3699 (.A(net3698),
    .X(net3699));
 sky130_fd_sc_hd__buf_1 place3582 (.A(_09100_),
    .X(net3582));
 sky130_fd_sc_hd__clkbuf_2 place3688 (.A(_09785_),
    .X(net3688));
 sky130_fd_sc_hd__clkbuf_2 place3685 (.A(_09935_),
    .X(net3685));
 sky130_fd_sc_hd__buf_1 place3684 (.A(_10057_),
    .X(net3684));
 sky130_fd_sc_hd__buf_1 place3683 (.A(_10131_),
    .X(net3683));
 sky130_fd_sc_hd__buf_8 rebuffer26 (.A(_08239_),
    .X(net281));
 sky130_fd_sc_hd__buf_1 place3584 (.A(_08631_),
    .X(net3584));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3586 (.A(_10547_),
    .X(net3586));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3690 (.A(_09721_),
    .X(net3690));
 sky130_fd_sc_hd__buf_12 place3676 (.A(_10332_),
    .X(net3676));
 sky130_fd_sc_hd__buf_1 place3675 (.A(_10415_),
    .X(net3675));
 sky130_fd_sc_hd__buf_1 place3673 (.A(_10541_),
    .X(net3673));
 sky130_fd_sc_hd__buf_1 place3679 (.A(net3677),
    .X(net3679));
 sky130_fd_sc_hd__buf_1 place3670 (.A(_02225_),
    .X(net3670));
 sky130_fd_sc_hd__buf_12 place3666 (.A(_08192_),
    .X(net3666));
 sky130_fd_sc_hd__buf_12 place3662 (.A(_12396_),
    .X(net3662));
 sky130_fd_sc_hd__buf_12 place3721 (.A(net293),
    .X(net3721));
 sky130_fd_sc_hd__clkbuf_2 place3661 (.A(net397),
    .X(net3661));
 sky130_fd_sc_hd__buf_1 place3807 (.A(net311),
    .X(net3807));
 sky130_fd_sc_hd__buf_12 place3795 (.A(net264),
    .X(net3795));
 sky130_fd_sc_hd__buf_12 place3803 (.A(_07983_),
    .X(net3803));
 sky130_fd_sc_hd__buf_8 place3800 (.A(net277),
    .X(net3800));
 sky130_fd_sc_hd__buf_6 place3657 (.A(_01689_),
    .X(net3657));
 sky130_fd_sc_hd__buf_1 place3654 (.A(net447),
    .X(net3654));
 sky130_fd_sc_hd__buf_12 place3861 (.A(net3860),
    .X(net3861));
 sky130_fd_sc_hd__buf_16 place3867 (.A(net3859),
    .X(net3867));
 sky130_fd_sc_hd__buf_12 place3866 (.A(net359),
    .X(net3866));
 sky130_fd_sc_hd__buf_1 place3640 (.A(_01794_),
    .X(net3640));
 sky130_fd_sc_hd__buf_12 place3639 (.A(_01843_),
    .X(net3639));
 sky130_fd_sc_hd__buf_6 place3645 (.A(_01771_),
    .X(net3645));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3648 (.A(_01758_),
    .X(net3648));
 sky130_fd_sc_hd__buf_12 place3895 (.A(net343),
    .X(net3895));
 sky130_fd_sc_hd__buf_1 place3636 (.A(_02318_),
    .X(net3636));
 sky130_fd_sc_hd__buf_2 place3894 (.A(net3893),
    .X(net3894));
 sky130_fd_sc_hd__buf_12 place3958 (.A(net3957),
    .X(net3958));
 sky130_fd_sc_hd__buf_12 place3893 (.A(net343),
    .X(net3893));
 sky130_fd_sc_hd__buf_1 place3892 (.A(net341),
    .X(net3892));
 sky130_fd_sc_hd__buf_2 place3881 (.A(net341),
    .X(net3881));
 sky130_fd_sc_hd__buf_12 place3629 (.A(_03307_),
    .X(net3629));
 sky130_fd_sc_hd__buf_1 place3628 (.A(net3627),
    .X(net3628));
 sky130_fd_sc_hd__buf_1 place3613 (.A(_09454_),
    .X(net3613));
 sky130_fd_sc_hd__buf_1 place3607 (.A(_01823_),
    .X(net3607));
 sky130_fd_sc_hd__buf_1 place3605 (.A(_01858_),
    .X(net3605));
 sky130_fd_sc_hd__buf_1 place3604 (.A(_01894_),
    .X(net3604));
 sky130_fd_sc_hd__buf_12 place3603 (.A(_02009_),
    .X(net3603));
 sky130_fd_sc_hd__buf_1 place3891 (.A(net343),
    .X(net3891));
 sky130_fd_sc_hd__clkbuf_2 place3890 (.A(net3888),
    .X(net3890));
 sky130_fd_sc_hd__buf_12 place3889 (.A(net3888),
    .X(net3889));
 sky130_fd_sc_hd__buf_1 place3592 (.A(_09107_),
    .X(net3592));
 sky130_fd_sc_hd__buf_1 place3593 (.A(_08954_),
    .X(net3593));
 sky130_fd_sc_hd__buf_12 place3917 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .X(net3917));
 sky130_fd_sc_hd__buf_1 place3589 (.A(_09371_),
    .X(net3589));
 sky130_fd_sc_hd__buf_1 place3590 (.A(_09310_),
    .X(net3590));
 sky130_fd_sc_hd__buf_1 place3587 (.A(_10427_),
    .X(net3587));
 sky130_fd_sc_hd__buf_16 place3930 (.A(net3929),
    .X(net3930));
 sky130_fd_sc_hd__buf_12 place3936 (.A(net3935),
    .X(net3936));
 sky130_fd_sc_hd__buf_12 place3962 (.A(net3961),
    .X(net3962));
 sky130_fd_sc_hd__buf_12 place3956 (.A(net3954),
    .X(net3956));
 sky130_fd_sc_hd__buf_12 place3961 (.A(net3960),
    .X(net3961));
 sky130_fd_sc_hd__buf_12 place3960 (.A(net148),
    .X(net3960));
 sky130_fd_sc_hd__buf_12 place3957 (.A(net148),
    .X(net3957));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3585 (.A(_01806_),
    .X(net3585));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3583 (.A(net484),
    .X(net3583));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3591 (.A(_09189_),
    .X(net3591));
 sky130_fd_sc_hd__buf_1 place3579 (.A(_01921_),
    .X(net3579));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__buf_2 place3874 (.A(net3873),
    .X(net3874));
 sky130_fd_sc_hd__buf_12 place3601 (.A(_08204_),
    .X(net3601));
 sky130_fd_sc_hd__buf_1 place3600 (.A(_08313_),
    .X(net3600));
 sky130_fd_sc_hd__buf_16 place3929 (.A(net3917),
    .X(net3929));
 sky130_fd_sc_hd__buf_1 place3599 (.A(_08410_),
    .X(net3599));
 sky130_fd_sc_hd__buf_8 place3597 (.A(_08545_),
    .X(net3597));
 sky130_fd_sc_hd__buf_1 place3595 (.A(net308),
    .X(net3595));
 sky130_fd_sc_hd__buf_12 place3920 (.A(net378),
    .X(net3920));
 sky130_fd_sc_hd__buf_12 place3594 (.A(_08709_),
    .X(net3594));
 sky130_fd_sc_hd__buf_12 place3973 (.A(net148),
    .X(net3973));
 sky130_fd_sc_hd__buf_1 place3596 (.A(_08621_),
    .X(net3596));
 sky130_fd_sc_hd__buf_12 place3598 (.A(net288),
    .X(net3598));
 sky130_fd_sc_hd__buf_12 place3888 (.A(net343),
    .X(net3888));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3602 (.A(_02122_),
    .X(net3602));
 sky130_fd_sc_hd__buf_12 place3972 (.A(net3971),
    .X(net3972));
 sky130_fd_sc_hd__buf_12 place3578 (.A(_02037_),
    .X(net3578));
 sky130_fd_sc_hd__buf_12 place3875 (.A(net3873),
    .X(net3875));
 sky130_fd_sc_hd__buf_12 place3577 (.A(_03691_),
    .X(net3577));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3609 (.A(_12418_),
    .X(net3609));
 sky130_fd_sc_hd__buf_1 place3574 (.A(_10719_),
    .X(net3574));
 sky130_fd_sc_hd__buf_1 place3572 (.A(_01922_),
    .X(net3572));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3573 (.A(_12170_),
    .X(net3573));
 sky130_fd_sc_hd__buf_1 place3570 (.A(_04051_),
    .X(net3570));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3568 (.A(_09112_),
    .X(net3568));
 sky130_fd_sc_hd__buf_1 place3565 (.A(_11309_),
    .X(net3565));
 sky130_fd_sc_hd__buf_1 place3563 (.A(_12174_),
    .X(net3563));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3560 (.A(_02013_),
    .X(net3560));
 sky130_fd_sc_hd__buf_12 place3559 (.A(_02016_),
    .X(net3559));
 sky130_fd_sc_hd__buf_1 place3557 (.A(_02171_),
    .X(net3557));
 sky130_fd_sc_hd__buf_1 place3552 (.A(_10604_),
    .X(net3552));
 sky130_fd_sc_hd__buf_1 place3551 (.A(_10607_),
    .X(net3551));
 sky130_fd_sc_hd__buf_12 place3550 (.A(_10615_),
    .X(net3550));
 sky130_fd_sc_hd__buf_1 place3549 (.A(net171),
    .X(net3549));
 sky130_fd_sc_hd__buf_1 place3547 (.A(_11059_),
    .X(net3547));
 sky130_fd_sc_hd__buf_1 place3546 (.A(_11070_),
    .X(net3546));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3543 (.A(_02278_),
    .X(net3543));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3537 (.A(net176),
    .X(net3537));
 sky130_fd_sc_hd__buf_6 place3533 (.A(_10710_),
    .X(net3533));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3530 (.A(net178),
    .X(net3530));
 sky130_fd_sc_hd__buf_12 place3529 (.A(_08815_),
    .X(net3529));
 sky130_fd_sc_hd__buf_1 place3522 (.A(_01997_),
    .X(net3522));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3520 (.A(net180),
    .X(net3520));
 sky130_fd_sc_hd__buf_12 place3534 (.A(net3533),
    .X(net3534));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3518 (.A(_02382_),
    .X(net3518));
 sky130_fd_sc_hd__buf_1 place3517 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .X(net3517));
 sky130_fd_sc_hd__buf_1 place3516 (.A(net152),
    .X(net3516));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3509 (.A(_02809_),
    .X(net3509));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3508 (.A(_02934_),
    .X(net3508));
 sky130_fd_sc_hd__buf_12 place3507 (.A(net156),
    .X(net3507));
 sky130_fd_sc_hd__buf_12 place3503 (.A(net163),
    .X(net3503));
 sky130_fd_sc_hd__buf_12 place3501 (.A(_10988_),
    .X(net3501));
 sky130_fd_sc_hd__buf_1 place3511 (.A(_09810_),
    .X(net3511));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3610 (.A(_12181_),
    .X(net3610));
 sky130_fd_sc_hd__buf_1 place3606 (.A(_01857_),
    .X(net3606));
 sky130_fd_sc_hd__buf_12 place3497 (.A(_09675_),
    .X(net3497));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3495 (.A(net166),
    .X(net3495));
 sky130_fd_sc_hd__buf_1 place3513 (.A(net155),
    .X(net3513));
 sky130_fd_sc_hd__buf_1 place3608 (.A(_01723_),
    .X(net3608));
 sky130_fd_sc_hd__buf_1 place3642 (.A(_01775_),
    .X(net3642));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3490 (.A(_11887_),
    .X(net3490));
 sky130_fd_sc_hd__buf_1 place3488 (.A(_03514_),
    .X(net3488));
 sky130_fd_sc_hd__bufbuf_16 place3486 (.A(_10242_),
    .X(net3486));
 sky130_fd_sc_hd__buf_1 place3485 (.A(_10372_),
    .X(net3485));
 sky130_fd_sc_hd__buf_12 place3484 (.A(_11147_),
    .X(net3484));
 sky130_fd_sc_hd__buf_1 place3483 (.A(_11441_),
    .X(net3483));
 sky130_fd_sc_hd__buf_1 place3482 (.A(_11476_),
    .X(net3482));
 sky130_fd_sc_hd__buf_1 place3481 (.A(_11490_),
    .X(net3481));
 sky130_fd_sc_hd__buf_8 place3536 (.A(net175),
    .X(net3536));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__buf_1 rebuffer154 (.A(net158),
    .X(net420));
 sky130_fd_sc_hd__buf_12 place3469 (.A(_01655_),
    .X(net3469));
 sky130_fd_sc_hd__buf_1 place3467 (.A(_04010_),
    .X(net3467));
 sky130_fd_sc_hd__buf_1 place3456 (.A(_05039_),
    .X(net3456));
 sky130_fd_sc_hd__buf_1 place3455 (.A(_05122_),
    .X(net3455));
 sky130_fd_sc_hd__buf_1 place3454 (.A(_07622_),
    .X(net3454));
 sky130_fd_sc_hd__buf_12 place3457 (.A(_04706_),
    .X(net3457));
 sky130_fd_sc_hd__buf_1 place3452 (.A(_04378_),
    .X(net3452));
 sky130_fd_sc_hd__buf_12 place3453 (.A(_02724_),
    .X(net3453));
 sky130_fd_sc_hd__buf_2 place3615 (.A(_08947_),
    .X(net3615));
 sky130_fd_sc_hd__buf_1 place3612 (.A(_10536_),
    .X(net3612));
 sky130_fd_sc_hd__buf_1 place3614 (.A(_09063_),
    .X(net3614));
 sky130_fd_sc_hd__buf_8 place3641 (.A(_01775_),
    .X(net3641));
 sky130_fd_sc_hd__buf_1 place3616 (.A(_08919_),
    .X(net3616));
 sky130_fd_sc_hd__buf_1 place3634 (.A(_02583_),
    .X(net3634));
 sky130_fd_sc_hd__buf_1 place3618 (.A(_08845_),
    .X(net3618));
 sky130_fd_sc_hd__buf_12 place3619 (.A(_08629_),
    .X(net3619));
 sky130_fd_sc_hd__buf_12 place3620 (.A(_08620_),
    .X(net3620));
 sky130_fd_sc_hd__buf_12 place3621 (.A(_08581_),
    .X(net3621));
 sky130_fd_sc_hd__buf_1 place3622 (.A(_08490_),
    .X(net3622));
 sky130_fd_sc_hd__buf_12 place3623 (.A(_08400_),
    .X(net3623));
 sky130_fd_sc_hd__buf_12 place3624 (.A(net290),
    .X(net3624));
 sky130_fd_sc_hd__buf_1 place3625 (.A(_08241_),
    .X(net3625));
 sky130_fd_sc_hd__buf_12 place3626 (.A(net300),
    .X(net3626));
 sky130_fd_sc_hd__buf_12 place3627 (.A(_03308_),
    .X(net3627));
 sky130_fd_sc_hd__buf_1 place3451 (.A(_04483_),
    .X(net3451));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net3762));
 sky130_fd_sc_hd__buf_12 place3631 (.A(_03058_),
    .X(net3631));
 sky130_fd_sc_hd__buf_1 place3632 (.A(_02784_),
    .X(net3632));
 sky130_fd_sc_hd__buf_1 place3450 (.A(_04731_),
    .X(net3450));
 sky130_fd_sc_hd__buf_1 place3544 (.A(_01995_),
    .X(net3544));
 sky130_fd_sc_hd__buf_12 place3635 (.A(_02324_),
    .X(net3635));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3545 (.A(_12178_),
    .X(net3545));
 sky130_fd_sc_hd__buf_1 place3651 (.A(_01711_),
    .X(net3651));
 sky130_fd_sc_hd__buf_1 place3652 (.A(_01705_),
    .X(net3652));
 sky130_fd_sc_hd__buf_1 place3653 (.A(_01705_),
    .X(net3653));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3637 (.A(_02236_),
    .X(net3637));
 sky130_fd_sc_hd__buf_12 place3655 (.A(net448),
    .X(net3655));
 sky130_fd_sc_hd__clkbuf_2 place3722 (.A(net3721),
    .X(net3722));
 sky130_fd_sc_hd__buf_12 place3638 (.A(_01867_),
    .X(net3638));
 sky130_fd_sc_hd__buf_12 place3443 (.A(net3440),
    .X(net3443));
 sky130_fd_sc_hd__buf_1 place3822 (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .X(net3822));
 sky130_fd_sc_hd__buf_1 place3946 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .X(net3946));
 sky130_fd_sc_hd__buf_1 place3856 (.A(net3854),
    .X(net3856));
 sky130_fd_sc_hd__buf_1 place3748 (.A(net321),
    .X(net3748));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3855 (.A(net3854),
    .X(net3855));
 sky130_fd_sc_hd__buf_12 place3845 (.A(net3844),
    .X(net3845));
 sky130_fd_sc_hd__buf_1 place3644 (.A(_01771_),
    .X(net3644));
 sky130_fd_sc_hd__buf_12 place3865 (.A(net3864),
    .X(net3865));
 sky130_fd_sc_hd__buf_1 place3944 (.A(net298),
    .X(net3944));
 sky130_fd_sc_hd__buf_1 place3824 (.A(\cs_registers_i.pc_id_i[28] ),
    .X(net3824));
 sky130_fd_sc_hd__buf_1 place3832 (.A(net286),
    .X(net3832));
 sky130_fd_sc_hd__buf_8 place3919 (.A(net346),
    .X(net3919));
 sky130_fd_sc_hd__clkbuf_2 place3646 (.A(_01765_),
    .X(net3646));
 sky130_fd_sc_hd__buf_12 place3918 (.A(net346),
    .X(net3918));
 sky130_fd_sc_hd__buf_12 place3847 (.A(net3844),
    .X(net3847));
 sky130_fd_sc_hd__buf_1 place3649 (.A(_01758_),
    .X(net3649));
 sky130_fd_sc_hd__buf_1 place3647 (.A(_01759_),
    .X(net3647));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__buf_1 place3650 (.A(net446),
    .X(net3650));
 sky130_fd_sc_hd__buf_12 place3928 (.A(net3927),
    .X(net3928));
 sky130_fd_sc_hd__buf_12 place3899 (.A(net349),
    .X(net3899));
 sky130_fd_sc_hd__buf_8 place3925 (.A(net3917),
    .X(net3925));
 sky130_fd_sc_hd__buf_1 place3943 (.A(net298),
    .X(net3943));
 sky130_fd_sc_hd__buf_16 place3924 (.A(net3922),
    .X(net3924));
 sky130_fd_sc_hd__buf_12 place3858 (.A(net360),
    .X(net3858));
 sky130_fd_sc_hd__buf_12 place3923 (.A(net3922),
    .X(net3923));
 sky130_fd_sc_hd__buf_1 place3805 (.A(net312),
    .X(net3805));
 sky130_fd_sc_hd__buf_12 place3898 (.A(net349),
    .X(net3898));
 sky130_fd_sc_hd__buf_16 place3927 (.A(net3917),
    .X(net3927));
 sky130_fd_sc_hd__buf_12 place3910 (.A(net3908),
    .X(net3910));
 sky130_fd_sc_hd__buf_1 place3897 (.A(net349),
    .X(net3897));
 sky130_fd_sc_hd__buf_12 place3911 (.A(net3908),
    .X(net3911));
 sky130_fd_sc_hd__buf_12 place3971 (.A(net148),
    .X(net3971));
 sky130_fd_sc_hd__buf_12 place3663 (.A(net3662),
    .X(net3663));
 sky130_fd_sc_hd__buf_12 place3979 (.A(net3974),
    .X(net3979));
 sky130_fd_sc_hd__buf_12 place3976 (.A(net3975),
    .X(net3976));
 sky130_fd_sc_hd__buf_12 place3975 (.A(net3974),
    .X(net3975));
 sky130_fd_sc_hd__buf_12 place3974 (.A(net148),
    .X(net3974));
 sky130_fd_sc_hd__buf_1 place3656 (.A(_01690_),
    .X(net3656));
 sky130_fd_sc_hd__buf_1 place3916 (.A(net3913),
    .X(net3916));
 sky130_fd_sc_hd__buf_1 place3887 (.A(net341),
    .X(net3887));
 sky130_fd_sc_hd__buf_8 place3864 (.A(net414),
    .X(net3864));
 sky130_fd_sc_hd__buf_12 place3863 (.A(net3860),
    .X(net3863));
 sky130_fd_sc_hd__buf_1 rebuffer123 (.A(net3917),
    .X(net378));
 sky130_fd_sc_hd__buf_1 place3659 (.A(_01683_),
    .X(net3659));
 sky130_fd_sc_hd__buf_12 place3658 (.A(net442),
    .X(net3658));
 sky130_fd_sc_hd__buf_6 place3860 (.A(net3859),
    .X(net3860));
 sky130_fd_sc_hd__buf_12 place3844 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .X(net3844));
 sky130_fd_sc_hd__buf_12 place3854 (.A(net256),
    .X(net3854));
 sky130_fd_sc_hd__buf_1 place3842 (.A(\id_stage_i.controller_i.instr_i[26] ),
    .X(net3842));
 sky130_fd_sc_hd__buf_1 place3660 (.A(net397),
    .X(net3660));
 sky130_fd_sc_hd__buf_1 place3841 (.A(net348),
    .X(net3841));
 sky130_fd_sc_hd__buf_1 place3840 (.A(net367),
    .X(net3840));
 sky130_fd_sc_hd__buf_1 place3843 (.A(\id_stage_i.controller_i.instr_i[25] ),
    .X(net3843));
 sky130_fd_sc_hd__buf_1 place3836 (.A(\id_stage_i.controller_i.instr_i[31] ),
    .X(net3836));
 sky130_fd_sc_hd__buf_1 place3711 (.A(net3710),
    .X(net3711));
 sky130_fd_sc_hd__buf_12 place3839 (.A(\id_stage_i.controller_i.instr_i[29] ),
    .X(net3839));
 sky130_fd_sc_hd__buf_1 place3834 (.A(net325),
    .X(net3834));
 sky130_fd_sc_hd__buf_1 place3835 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net3835));
 sky130_fd_sc_hd__buf_1 place3680 (.A(_10229_),
    .X(net3680));
 sky130_fd_sc_hd__buf_1 place3664 (.A(net369),
    .X(net3664));
 sky130_fd_sc_hd__buf_1 place3825 (.A(\cs_registers_i.pc_id_i[27] ),
    .X(net3825));
 sky130_fd_sc_hd__buf_1 place3821 (.A(_07845_),
    .X(net3821));
 sky130_fd_sc_hd__buf_8 place3852 (.A(net256),
    .X(net3852));
 sky130_fd_sc_hd__buf_1 place3838 (.A(\id_stage_i.controller_i.instr_i[2] ),
    .X(net3838));
 sky130_fd_sc_hd__buf_1 place3827 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .X(net3827));
 sky130_fd_sc_hd__buf_12 place3665 (.A(_08202_),
    .X(net3665));
 sky130_fd_sc_hd__buf_12 place3859 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .X(net3859));
 sky130_fd_sc_hd__buf_1 place3671 (.A(_01687_),
    .X(net3671));
 sky130_fd_sc_hd__buf_1 place3667 (.A(_07912_),
    .X(net3667));
 sky130_fd_sc_hd__buf_12 place3809 (.A(_07969_),
    .X(net3809));
 sky130_fd_sc_hd__buf_12 place3668 (.A(_03681_),
    .X(net3668));
 sky130_fd_sc_hd__buf_2 place3710 (.A(net3709),
    .X(net3710));
 sky130_fd_sc_hd__buf_1 place3691 (.A(_09704_),
    .X(net3691));
 sky130_fd_sc_hd__buf_1 place3678 (.A(net3677),
    .X(net3678));
 sky130_fd_sc_hd__buf_12 place3804 (.A(net313),
    .X(net3804));
 sky130_fd_sc_hd__buf_12 place3802 (.A(_07983_),
    .X(net3802));
 sky130_fd_sc_hd__buf_12 place3810 (.A(_07962_),
    .X(net3810));
 sky130_fd_sc_hd__buf_1 place3672 (.A(_13078_),
    .X(net3672));
 sky130_fd_sc_hd__buf_1 place3833 (.A(net325),
    .X(net3833));
 sky130_fd_sc_hd__buf_12 place3677 (.A(_10265_),
    .X(net3677));
 sky130_fd_sc_hd__buf_12 place3681 (.A(_10199_),
    .X(net3681));
 sky130_fd_sc_hd__buf_1 place3682 (.A(_10157_),
    .X(net3682));
 sky130_fd_sc_hd__buf_1 place3823 (.A(\cs_registers_i.pc_id_i[8] ),
    .X(net3823));
 sky130_fd_sc_hd__clkbuf_2 place3819 (.A(_07856_),
    .X(net3819));
 sky130_fd_sc_hd__buf_2 place3799 (.A(_07993_),
    .X(net3799));
 sky130_fd_sc_hd__buf_1 place3831 (.A(net286),
    .X(net3831));
 sky130_fd_sc_hd__buf_1 place3686 (.A(_09863_),
    .X(net3686));
 sky130_fd_sc_hd__buf_12 place3798 (.A(_07993_),
    .X(net3798));
 sky130_fd_sc_hd__buf_1 place3797 (.A(_08056_),
    .X(net3797));
 sky130_fd_sc_hd__buf_1 place3689 (.A(_09760_),
    .X(net3689));
 sky130_fd_sc_hd__buf_2 place3692 (.A(_09620_),
    .X(net3692));
 sky130_fd_sc_hd__buf_2 place3796 (.A(_08135_),
    .X(net3796));
 sky130_fd_sc_hd__buf_2 place3791 (.A(_08147_),
    .X(net3791));
 sky130_fd_sc_hd__buf_1 place3789 (.A(net3788),
    .X(net3789));
 sky130_fd_sc_hd__buf_1 place3786 (.A(_08171_),
    .X(net3786));
 sky130_fd_sc_hd__buf_12 place3784 (.A(_08258_),
    .X(net3784));
 sky130_fd_sc_hd__buf_12 place3693 (.A(net310),
    .X(net3693));
 sky130_fd_sc_hd__buf_12 place3698 (.A(_09181_),
    .X(net3698));
 sky130_fd_sc_hd__buf_12 place3788 (.A(_08158_),
    .X(net3788));
 sky130_fd_sc_hd__buf_12 place3696 (.A(_09335_),
    .X(net3696));
 sky130_fd_sc_hd__buf_1 place3703 (.A(net3702),
    .X(net3703));
 sky130_fd_sc_hd__buf_12 place3697 (.A(_09302_),
    .X(net3697));
 sky130_fd_sc_hd__buf_1 place3829 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .X(net3829));
 sky130_fd_sc_hd__buf_8 place3709 (.A(_08616_),
    .X(net3709));
 sky130_fd_sc_hd__buf_12 place3785 (.A(_08181_),
    .X(net3785));
 sky130_fd_sc_hd__buf_1 place3701 (.A(_09062_),
    .X(net3701));
 sky130_fd_sc_hd__buf_1 place3783 (.A(_08261_),
    .X(net3783));
 sky130_fd_sc_hd__buf_1 place3782 (.A(_08266_),
    .X(net3782));
 sky130_fd_sc_hd__buf_12 place3702 (.A(_08985_),
    .X(net3702));
 sky130_fd_sc_hd__buf_1 place3704 (.A(_08939_),
    .X(net3704));
 sky130_fd_sc_hd__buf_12 place3781 (.A(_08279_),
    .X(net3781));
 sky130_fd_sc_hd__buf_2 place3706 (.A(net340),
    .X(net3706));
 sky130_fd_sc_hd__buf_12 place3707 (.A(_08733_),
    .X(net3707));
 sky130_fd_sc_hd__buf_12 place3778 (.A(net370),
    .X(net3778));
 sky130_fd_sc_hd__buf_1 place3708 (.A(_08703_),
    .X(net3708));
 sky130_fd_sc_hd__buf_12 place3712 (.A(_08574_),
    .X(net3712));
 sky130_fd_sc_hd__buf_1 place3714 (.A(net3713),
    .X(net3714));
 sky130_fd_sc_hd__buf_4 place3715 (.A(_08488_),
    .X(net3715));
 sky130_fd_sc_hd__buf_1 place3720 (.A(net293),
    .X(net3720));
 sky130_fd_sc_hd__buf_1 place3717 (.A(net3716),
    .X(net3717));
 sky130_fd_sc_hd__buf_8 place3769 (.A(_08522_),
    .X(net3769));
 sky130_fd_sc_hd__buf_12 place3719 (.A(_08346_),
    .X(net3719));
 sky130_fd_sc_hd__buf_12 place3716 (.A(_08394_),
    .X(net3716));
 sky130_fd_sc_hd__buf_8 place3816 (.A(net345),
    .X(net3816));
 sky130_fd_sc_hd__buf_1 place3718 (.A(_08348_),
    .X(net3718));
 sky130_fd_sc_hd__buf_1 place3775 (.A(net260),
    .X(net3775));
 sky130_fd_sc_hd__buf_1 place3724 (.A(net435),
    .X(net3724));
 sky130_fd_sc_hd__buf_2 place3749 (.A(_08194_),
    .X(net3749));
 sky130_fd_sc_hd__buf_8 place3726 (.A(net416),
    .X(net3726));
 sky130_fd_sc_hd__buf_6 place3727 (.A(_07999_),
    .X(net3727));
 sky130_fd_sc_hd__buf_1 place3734 (.A(_10690_),
    .X(net3734));
 sky130_fd_sc_hd__buf_1 place3729 (.A(_07045_),
    .X(net3729));
 sky130_fd_sc_hd__buf_12 place3752 (.A(_07960_),
    .X(net3752));
 sky130_fd_sc_hd__buf_12 place3738 (.A(_08406_),
    .X(net3738));
 sky130_fd_sc_hd__buf_12 place3739 (.A(_08316_),
    .X(net3739));
 sky130_fd_sc_hd__buf_1 place3740 (.A(_07894_),
    .X(net3740));
 sky130_fd_sc_hd__buf_12 place3742 (.A(_10777_),
    .X(net3742));
 sky130_fd_sc_hd__buf_1 place3743 (.A(net321),
    .X(net3743));
 sky130_fd_sc_hd__buf_1 place3761 (.A(_01677_),
    .X(net3761));
 sky130_fd_sc_hd__buf_12 place3757 (.A(_01708_),
    .X(net3757));
 sky130_fd_sc_hd__buf_1 place3820 (.A(_07850_),
    .X(net3820));
 sky130_fd_sc_hd__buf_8 place3768 (.A(_08531_),
    .X(net3768));
 sky130_fd_sc_hd__buf_8 place3770 (.A(_08391_),
    .X(net3770));
 sky130_fd_sc_hd__buf_12 place3755 (.A(_07857_),
    .X(net3755));
 sky130_fd_sc_hd__buf_12 place3754 (.A(_07872_),
    .X(net3754));
 sky130_fd_sc_hd__buf_8 place3772 (.A(_08299_),
    .X(net3772));
 sky130_fd_sc_hd__buf_1 place3771 (.A(_08374_),
    .X(net3771));
 sky130_fd_sc_hd__buf_12 place3794 (.A(net266),
    .X(net3794));
 sky130_fd_sc_hd__buf_1 place3828 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .X(net3828));
 sky130_fd_sc_hd__buf_1 place3790 (.A(_08147_),
    .X(net3790));
 sky130_fd_sc_hd__buf_12 place3793 (.A(net265),
    .X(net3793));
 sky130_fd_sc_hd__buf_12 place3806 (.A(net311),
    .X(net3806));
 sky130_fd_sc_hd__buf_12 place3801 (.A(net278),
    .X(net3801));
 sky130_fd_sc_hd__buf_12 place3808 (.A(_07969_),
    .X(net3808));
 sky130_fd_sc_hd__buf_12 place3811 (.A(_07962_),
    .X(net3811));
 sky130_fd_sc_hd__buf_4 place3815 (.A(net395),
    .X(net3815));
 sky130_fd_sc_hd__clkbuf_2 place3812 (.A(_07955_),
    .X(net3812));
 sky130_fd_sc_hd__buf_8 place3814 (.A(net364),
    .X(net3814));
 sky130_fd_sc_hd__buf_6 place3813 (.A(net365),
    .X(net3813));
 sky130_fd_sc_hd__buf_12 place3849 (.A(net3848),
    .X(net3849));
 sky130_fd_sc_hd__buf_1 place3818 (.A(_07885_),
    .X(net3818));
 sky130_fd_sc_hd__buf_12 place3848 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .X(net3848));
 sky130_fd_sc_hd__buf_8 place3830 (.A(\id_stage_i.controller_i.instr_i[6] ),
    .X(net3830));
 sky130_fd_sc_hd__buf_1 place3837 (.A(net355),
    .X(net3837));
 sky130_fd_sc_hd__buf_12 place3915 (.A(net3914),
    .X(net3915));
 sky130_fd_sc_hd__buf_12 place3885 (.A(net3884),
    .X(net3885));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__buf_12 place3882 (.A(net343),
    .X(net3882));
 sky130_fd_sc_hd__buf_1 place3942 (.A(net298),
    .X(net3942));
 sky130_fd_sc_hd__buf_1 place3938 (.A(net356),
    .X(net3938));
 sky130_fd_sc_hd__buf_12 place3901 (.A(net3900),
    .X(net3901));
 sky130_fd_sc_hd__buf_12 place3965 (.A(net3964),
    .X(net3965));
 sky130_fd_sc_hd__buf_16 place3926 (.A(net3917),
    .X(net3926));
 sky130_fd_sc_hd__buf_12 place3846 (.A(net3844),
    .X(net3846));
 sky130_fd_sc_hd__buf_12 place3959 (.A(net148),
    .X(net3959));
 sky130_fd_sc_hd__buf_12 place3935 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .X(net3935));
 sky130_fd_sc_hd__buf_12 place3939 (.A(net357),
    .X(net3939));
 sky130_fd_sc_hd__clkbuf_4 place3909 (.A(net3908),
    .X(net3909));
 sky130_fd_sc_hd__buf_1 place3905 (.A(net3902),
    .X(net3905));
 sky130_fd_sc_hd__buf_12 place3904 (.A(net3903),
    .X(net3904));
 sky130_fd_sc_hd__buf_12 place3902 (.A(net283),
    .X(net3902));
 sky130_fd_sc_hd__buf_12 place3908 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net3908));
 sky130_fd_sc_hd__buf_12 place3903 (.A(net3902),
    .X(net3903));
 sky130_fd_sc_hd__buf_1 place3941 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net3941));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__conb_1 _26833__6 (.LO(net255));
 sky130_fd_sc_hd__buf_12 place3968 (.A(net3967),
    .X(net3968));
 sky130_fd_sc_hd__conb_1 _26800__3 (.LO(net252));
 sky130_fd_sc_hd__conb_1 ibex_core_1 (.LO(net250));
 sky130_fd_sc_hd__buf_12 place3954 (.A(net148),
    .X(net3954));
 sky130_fd_sc_hd__buf_1 place3945 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .X(net3945));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_08275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_08275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_08437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_08437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net3803));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net3713));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net3713));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_08939_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_08939_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_09038_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_09730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_09903_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_10088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_10736_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_11398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_11726_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(boot_addr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(boot_addr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(boot_addr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(boot_addr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(boot_addr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(boot_addr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(data_rdata_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(fetch_enable_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(hart_id_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(hart_id_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(hart_id_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(irq_fast_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(irq_fast_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(irq_fast_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net3809));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net3802));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net3677));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net3682));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net3702));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net3702));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net3704));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net3793));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net3848));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_08167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net3929));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_10088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\cs_registers_i.csr_depc_o[25] ));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1134 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_900 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1137 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1082 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1080 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_962 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1134 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1080 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1194 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1100 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1052 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_954 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_962 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_962 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1142 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_924 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_983 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1020 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_954 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1187 ();
 assign alert_major_o = net250;
endmodule
