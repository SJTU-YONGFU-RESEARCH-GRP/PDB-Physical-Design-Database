module configurable_priority_encoder (valid,
    grant_index,
    request);
 output valid;
 output [2:0] grant_index;
 input [7:0] request;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12_ (.I(net2),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13_ (.I(net7),
    .ZN(_01_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14_ (.A1(_01_),
    .A2(net8),
    .B(net6),
    .ZN(_02_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15_ (.A1(net1),
    .A2(net5),
    .A3(net3),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16_ (.I(net1),
    .ZN(_04_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17_ (.A1(_04_),
    .A2(net4),
    .ZN(_05_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _18_ (.A1(net1),
    .A2(_00_),
    .B1(_02_),
    .B2(_03_),
    .C1(_05_),
    .C2(net3),
    .ZN(net9));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19_ (.A1(net4),
    .A2(net3),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20_ (.A1(net7),
    .A2(net8),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21_ (.A1(net6),
    .A2(net5),
    .A3(_07_),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22_ (.A1(_06_),
    .A2(_08_),
    .B(net1),
    .C(net2),
    .ZN(net10));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23_ (.A1(net6),
    .A2(net5),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24_ (.A1(_07_),
    .A2(_09_),
    .ZN(_10_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25_ (.A1(_04_),
    .A2(_00_),
    .A3(_06_),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26_ (.A1(_10_),
    .A2(_11_),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27_ (.A1(_07_),
    .A2(_09_),
    .A3(_11_),
    .ZN(net12));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_42 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_52 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input1 (.I(request[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(request[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input3 (.I(request[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(request[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(request[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(request[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(request[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(request[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net9),
    .Z(grant_index[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net10),
    .Z(grant_index[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net11),
    .Z(grant_index[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net12),
    .Z(valid));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_192 ();
endmodule
