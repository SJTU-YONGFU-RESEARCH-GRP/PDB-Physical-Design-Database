module sipo_register (clk,
    enable,
    parity_out,
    rst_n,
    serial_in,
    parallel_out);
 input clk;
 input enable;
 output parity_out;
 input rst_n;
 input serial_in;
 output [7:0] parallel_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X2 _36_ (.A(rst_n),
    .Z(_09_));
 CLKBUF_X3 _37_ (.A(enable),
    .Z(_10_));
 OAI21_X1 _38_ (.A(_09_),
    .B1(_10_),
    .B2(net10),
    .ZN(_11_));
 XNOR2_X1 _39_ (.A(net7),
    .B(net8),
    .ZN(_12_));
 XNOR2_X1 _40_ (.A(net5),
    .B(net6),
    .ZN(_13_));
 XNOR2_X1 _41_ (.A(_12_),
    .B(_13_),
    .ZN(_14_));
 XNOR2_X1 _42_ (.A(net3),
    .B(net4),
    .ZN(_15_));
 XNOR2_X1 _43_ (.A(net2),
    .B(net1),
    .ZN(_16_));
 XNOR2_X1 _44_ (.A(_15_),
    .B(_16_),
    .ZN(_17_));
 XNOR2_X1 _45_ (.A(_14_),
    .B(_17_),
    .ZN(_18_));
 AOI21_X1 _46_ (.A(_11_),
    .B1(_18_),
    .B2(_10_),
    .ZN(_00_));
 MUX2_X1 _47_ (.A(net2),
    .B(net1),
    .S(_10_),
    .Z(_19_));
 AND2_X1 _48_ (.A1(_09_),
    .A2(_19_),
    .ZN(_01_));
 MUX2_X1 _49_ (.A(net3),
    .B(net2),
    .S(_10_),
    .Z(_20_));
 AND2_X1 _50_ (.A1(_09_),
    .A2(_20_),
    .ZN(_02_));
 MUX2_X1 _51_ (.A(net4),
    .B(net3),
    .S(_10_),
    .Z(_21_));
 AND2_X1 _52_ (.A1(_09_),
    .A2(_21_),
    .ZN(_03_));
 MUX2_X1 _53_ (.A(net5),
    .B(net4),
    .S(_10_),
    .Z(_22_));
 AND2_X1 _54_ (.A1(_09_),
    .A2(_22_),
    .ZN(_04_));
 MUX2_X1 _55_ (.A(net6),
    .B(net5),
    .S(_10_),
    .Z(_23_));
 AND2_X1 _56_ (.A1(_09_),
    .A2(_23_),
    .ZN(_05_));
 MUX2_X1 _57_ (.A(net7),
    .B(net6),
    .S(_10_),
    .Z(_24_));
 AND2_X1 _58_ (.A1(_09_),
    .A2(_24_),
    .ZN(_06_));
 MUX2_X1 _59_ (.A(net8),
    .B(net7),
    .S(_10_),
    .Z(_25_));
 AND2_X1 _60_ (.A1(_09_),
    .A2(_25_),
    .ZN(_07_));
 MUX2_X1 _61_ (.A(net9),
    .B(net8),
    .S(_10_),
    .Z(_26_));
 AND2_X1 _62_ (.A1(_09_),
    .A2(_26_),
    .ZN(_08_));
 DFF_X1 \parity_bit$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net10),
    .QN(_35_));
 DFF_X1 \shift_reg[0]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net2),
    .QN(_34_));
 DFF_X1 \shift_reg[1]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net3),
    .QN(_33_));
 DFF_X1 \shift_reg[2]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_32_));
 DFF_X1 \shift_reg[3]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_31_));
 DFF_X1 \shift_reg[4]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net6),
    .QN(_30_));
 DFF_X1 \shift_reg[5]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net7),
    .QN(_29_));
 DFF_X1 \shift_reg[6]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net8),
    .QN(_28_));
 DFF_X1 \shift_reg[7]$_SDFFE_PN0P_  (.D(_08_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net9),
    .QN(_27_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_55 ();
 BUF_X1 input1 (.A(serial_in),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(parallel_out[0]));
 BUF_X1 output3 (.A(net3),
    .Z(parallel_out[1]));
 BUF_X1 output4 (.A(net4),
    .Z(parallel_out[2]));
 BUF_X1 output5 (.A(net5),
    .Z(parallel_out[3]));
 BUF_X1 output6 (.A(net6),
    .Z(parallel_out[4]));
 BUF_X1 output7 (.A(net7),
    .Z(parallel_out[5]));
 BUF_X1 output8 (.A(net8),
    .Z(parallel_out[6]));
 BUF_X1 output9 (.A(net9),
    .Z(parallel_out[7]));
 BUF_X1 output10 (.A(net10),
    .Z(parity_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X8 FILLER_0_92 ();
 FILLCELL_X4 FILLER_0_100 ();
 FILLCELL_X2 FILLER_0_104 ();
 FILLCELL_X8 FILLER_0_109 ();
 FILLCELL_X2 FILLER_0_117 ();
 FILLCELL_X32 FILLER_0_122 ();
 FILLCELL_X32 FILLER_0_154 ();
 FILLCELL_X16 FILLER_0_186 ();
 FILLCELL_X4 FILLER_0_202 ();
 FILLCELL_X2 FILLER_0_206 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X1 FILLER_1_81 ();
 FILLCELL_X2 FILLER_1_86 ();
 FILLCELL_X32 FILLER_1_105 ();
 FILLCELL_X32 FILLER_1_137 ();
 FILLCELL_X32 FILLER_1_169 ();
 FILLCELL_X4 FILLER_1_201 ();
 FILLCELL_X2 FILLER_1_205 ();
 FILLCELL_X1 FILLER_1_207 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_89 ();
 FILLCELL_X1 FILLER_2_95 ();
 FILLCELL_X32 FILLER_2_130 ();
 FILLCELL_X32 FILLER_2_162 ();
 FILLCELL_X8 FILLER_2_194 ();
 FILLCELL_X4 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_206 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X16 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_81 ();
 FILLCELL_X2 FILLER_3_85 ();
 FILLCELL_X1 FILLER_3_87 ();
 FILLCELL_X1 FILLER_3_95 ();
 FILLCELL_X1 FILLER_3_103 ();
 FILLCELL_X1 FILLER_3_110 ();
 FILLCELL_X1 FILLER_3_118 ();
 FILLCELL_X32 FILLER_3_123 ();
 FILLCELL_X32 FILLER_3_155 ();
 FILLCELL_X16 FILLER_3_187 ();
 FILLCELL_X4 FILLER_3_203 ();
 FILLCELL_X1 FILLER_3_207 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X16 FILLER_4_65 ();
 FILLCELL_X8 FILLER_4_81 ();
 FILLCELL_X4 FILLER_4_89 ();
 FILLCELL_X1 FILLER_4_93 ();
 FILLCELL_X32 FILLER_4_110 ();
 FILLCELL_X32 FILLER_4_142 ();
 FILLCELL_X32 FILLER_4_174 ();
 FILLCELL_X2 FILLER_4_206 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X8 FILLER_5_97 ();
 FILLCELL_X2 FILLER_5_105 ();
 FILLCELL_X1 FILLER_5_107 ();
 FILLCELL_X32 FILLER_5_116 ();
 FILLCELL_X32 FILLER_5_148 ();
 FILLCELL_X16 FILLER_5_180 ();
 FILLCELL_X8 FILLER_5_196 ();
 FILLCELL_X4 FILLER_5_204 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X8 FILLER_6_193 ();
 FILLCELL_X4 FILLER_6_201 ();
 FILLCELL_X2 FILLER_6_205 ();
 FILLCELL_X1 FILLER_6_207 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_81 ();
 FILLCELL_X2 FILLER_7_85 ();
 FILLCELL_X1 FILLER_7_87 ();
 FILLCELL_X8 FILLER_7_92 ();
 FILLCELL_X4 FILLER_7_100 ();
 FILLCELL_X2 FILLER_7_104 ();
 FILLCELL_X1 FILLER_7_106 ();
 FILLCELL_X32 FILLER_7_114 ();
 FILLCELL_X32 FILLER_7_146 ();
 FILLCELL_X16 FILLER_7_178 ();
 FILLCELL_X8 FILLER_7_194 ();
 FILLCELL_X4 FILLER_7_202 ();
 FILLCELL_X2 FILLER_7_206 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_81 ();
 FILLCELL_X1 FILLER_8_85 ();
 FILLCELL_X1 FILLER_8_103 ();
 FILLCELL_X32 FILLER_8_125 ();
 FILLCELL_X32 FILLER_8_157 ();
 FILLCELL_X16 FILLER_8_189 ();
 FILLCELL_X2 FILLER_8_205 ();
 FILLCELL_X1 FILLER_8_207 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X2 FILLER_9_81 ();
 FILLCELL_X8 FILLER_9_90 ();
 FILLCELL_X2 FILLER_9_98 ();
 FILLCELL_X1 FILLER_9_100 ();
 FILLCELL_X32 FILLER_9_106 ();
 FILLCELL_X32 FILLER_9_138 ();
 FILLCELL_X32 FILLER_9_170 ();
 FILLCELL_X4 FILLER_9_202 ();
 FILLCELL_X2 FILLER_9_206 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X8 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_172 ();
 FILLCELL_X4 FILLER_10_204 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X16 FILLER_11_65 ();
 FILLCELL_X1 FILLER_11_81 ();
 FILLCELL_X32 FILLER_11_99 ();
 FILLCELL_X32 FILLER_11_131 ();
 FILLCELL_X32 FILLER_11_163 ();
 FILLCELL_X8 FILLER_11_195 ();
 FILLCELL_X4 FILLER_11_203 ();
 FILLCELL_X1 FILLER_11_207 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X16 FILLER_12_65 ();
 FILLCELL_X1 FILLER_12_81 ();
 FILLCELL_X2 FILLER_12_93 ();
 FILLCELL_X32 FILLER_12_100 ();
 FILLCELL_X32 FILLER_12_132 ();
 FILLCELL_X32 FILLER_12_164 ();
 FILLCELL_X8 FILLER_12_196 ();
 FILLCELL_X4 FILLER_12_204 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_81 ();
 FILLCELL_X1 FILLER_13_105 ();
 FILLCELL_X32 FILLER_13_112 ();
 FILLCELL_X32 FILLER_13_144 ();
 FILLCELL_X32 FILLER_13_176 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X8 FILLER_14_65 ();
 FILLCELL_X4 FILLER_14_73 ();
 FILLCELL_X2 FILLER_14_77 ();
 FILLCELL_X1 FILLER_14_79 ();
 FILLCELL_X1 FILLER_14_88 ();
 FILLCELL_X4 FILLER_14_96 ();
 FILLCELL_X1 FILLER_14_100 ();
 FILLCELL_X4 FILLER_14_107 ();
 FILLCELL_X1 FILLER_14_111 ();
 FILLCELL_X2 FILLER_14_116 ();
 FILLCELL_X1 FILLER_14_118 ();
 FILLCELL_X32 FILLER_14_123 ();
 FILLCELL_X32 FILLER_14_155 ();
 FILLCELL_X16 FILLER_14_187 ();
 FILLCELL_X4 FILLER_14_203 ();
 FILLCELL_X1 FILLER_14_207 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_69 ();
 FILLCELL_X1 FILLER_15_71 ();
 FILLCELL_X2 FILLER_15_96 ();
 FILLCELL_X4 FILLER_15_104 ();
 FILLCELL_X1 FILLER_15_125 ();
 FILLCELL_X32 FILLER_15_131 ();
 FILLCELL_X32 FILLER_15_163 ();
 FILLCELL_X8 FILLER_15_195 ();
 FILLCELL_X4 FILLER_15_203 ();
 FILLCELL_X1 FILLER_15_207 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_9 ();
 FILLCELL_X1 FILLER_16_11 ();
 FILLCELL_X32 FILLER_16_15 ();
 FILLCELL_X32 FILLER_16_47 ();
 FILLCELL_X32 FILLER_16_79 ();
 FILLCELL_X32 FILLER_16_111 ();
 FILLCELL_X16 FILLER_16_143 ();
 FILLCELL_X8 FILLER_16_159 ();
 FILLCELL_X2 FILLER_16_167 ();
 FILLCELL_X1 FILLER_16_169 ();
 FILLCELL_X32 FILLER_16_173 ();
 FILLCELL_X2 FILLER_16_205 ();
 FILLCELL_X1 FILLER_16_207 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X8 FILLER_17_193 ();
 FILLCELL_X4 FILLER_17_201 ();
 FILLCELL_X2 FILLER_17_205 ();
 FILLCELL_X1 FILLER_17_207 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X8 FILLER_18_193 ();
 FILLCELL_X4 FILLER_18_201 ();
 FILLCELL_X2 FILLER_18_205 ();
 FILLCELL_X1 FILLER_18_207 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X8 FILLER_19_193 ();
 FILLCELL_X4 FILLER_19_201 ();
 FILLCELL_X2 FILLER_19_205 ();
 FILLCELL_X1 FILLER_19_207 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X8 FILLER_20_193 ();
 FILLCELL_X4 FILLER_20_201 ();
 FILLCELL_X2 FILLER_20_205 ();
 FILLCELL_X1 FILLER_20_207 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X8 FILLER_21_193 ();
 FILLCELL_X4 FILLER_21_201 ();
 FILLCELL_X2 FILLER_21_205 ();
 FILLCELL_X1 FILLER_21_207 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X8 FILLER_22_193 ();
 FILLCELL_X4 FILLER_22_201 ();
 FILLCELL_X2 FILLER_22_205 ();
 FILLCELL_X1 FILLER_22_207 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_193 ();
 FILLCELL_X4 FILLER_23_201 ();
 FILLCELL_X2 FILLER_23_205 ();
 FILLCELL_X1 FILLER_23_207 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X8 FILLER_24_193 ();
 FILLCELL_X4 FILLER_24_201 ();
 FILLCELL_X2 FILLER_24_205 ();
 FILLCELL_X1 FILLER_24_207 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X8 FILLER_25_193 ();
 FILLCELL_X4 FILLER_25_201 ();
 FILLCELL_X2 FILLER_25_205 ();
 FILLCELL_X1 FILLER_25_207 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X16 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_81 ();
 FILLCELL_X2 FILLER_26_85 ();
 FILLCELL_X32 FILLER_26_90 ();
 FILLCELL_X32 FILLER_26_122 ();
 FILLCELL_X32 FILLER_26_154 ();
 FILLCELL_X16 FILLER_26_186 ();
 FILLCELL_X4 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_206 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X4 FILLER_27_81 ();
 FILLCELL_X1 FILLER_27_85 ();
 FILLCELL_X2 FILLER_27_89 ();
 FILLCELL_X32 FILLER_27_94 ();
 FILLCELL_X32 FILLER_27_126 ();
 FILLCELL_X32 FILLER_27_158 ();
 FILLCELL_X16 FILLER_27_190 ();
 FILLCELL_X2 FILLER_27_206 ();
endmodule
