module circular_buffer_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    peek_en,
    rd_en,
    rst_n,
    wr_en,
    fifo_count,
    peek_addr,
    peek_data,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input peek_en;
 input rd_en;
 input rst_n;
 input wr_en;
 output [4:0] fifo_count;
 input [3:0] peek_addr;
 output [7:0] peek_data;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net42;

 sky130_fd_sc_hd__inv_1 _259_ (.A(net21),
    .Y(_245_));
 sky130_fd_sc_hd__nand3b_2 _260_ (.A_N(_257_),
    .B(_235_),
    .C(_238_),
    .Y(_037_));
 sky130_fd_sc_hd__a21oi_2 _261_ (.A1(_238_),
    .A2(_234_),
    .B1(_237_),
    .Y(_038_));
 sky130_fd_sc_hd__a21boi_2 _262_ (.A1(_037_),
    .A2(_038_),
    .B1_N(_233_),
    .Y(_039_));
 sky130_fd_sc_hd__and3b_1 _263_ (.A_N(_257_),
    .B(_235_),
    .C(_238_),
    .X(_040_));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(_238_),
    .A2(_234_),
    .B1(_237_),
    .X(_041_));
 sky130_fd_sc_hd__nor3_2 _265_ (.A(_233_),
    .B(_040_),
    .C(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _266_ (.A(_039_),
    .B(_042_),
    .Y(net23));
 sky130_fd_sc_hd__xor2_2 _267_ (.A(_238_),
    .B(_226_),
    .X(net22));
 sky130_fd_sc_hd__inv_1 _268_ (.A(_258_),
    .Y(net20));
 sky130_fd_sc_hd__a21o_1 _269_ (.A1(_238_),
    .A2(_226_),
    .B1(_237_),
    .X(_043_));
 sky130_fd_sc_hd__a21oi_2 _270_ (.A1(_233_),
    .A2(_043_),
    .B1(_232_),
    .Y(_044_));
 sky130_fd_sc_hd__xnor2_2 _271_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Y(_045_));
 sky130_fd_sc_hd__xnor2_4 _272_ (.A(_044_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__buf_4 _273_ (.A(_046_),
    .X(net24));
 sky130_fd_sc_hd__nor3_1 _274_ (.A(net20),
    .B(net21),
    .C(net22),
    .Y(_047_));
 sky130_fd_sc_hd__o21a_2 _275_ (.A1(_039_),
    .A2(_042_),
    .B1(_047_),
    .X(_048_));
 sky130_fd_sc_hd__and2_0 _276_ (.A(net24),
    .B(_048_),
    .X(net25));
 sky130_fd_sc_hd__o21ai_4 _277_ (.A1(_039_),
    .A2(_042_),
    .B1(_047_),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_1 _278_ (.A(net24),
    .B(_049_),
    .Y(net19));
 sky130_fd_sc_hd__and2_0 _279_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .X(_050_));
 sky130_fd_sc_hd__inv_1 _280_ (.A(net16),
    .Y(_051_));
 sky130_fd_sc_hd__a21oi_2 _281_ (.A1(_046_),
    .A2(_048_),
    .B1(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__and3_4 _282_ (.A(_250_),
    .B(_050_),
    .C(_052_),
    .X(_003_));
 sky130_fd_sc_hd__and3_4 _283_ (.A(_253_),
    .B(_050_),
    .C(_052_),
    .X(_004_));
 sky130_fd_sc_hd__and3_4 _284_ (.A(_251_),
    .B(_050_),
    .C(_052_),
    .X(_005_));
 sky130_fd_sc_hd__nand3_1 _285_ (.A(net16),
    .B(_255_),
    .C(_050_),
    .Y(_053_));
 sky130_fd_sc_hd__a21oi_4 _286_ (.A1(_046_),
    .A2(_048_),
    .B1(_053_),
    .Y(_006_));
 sky130_fd_sc_hd__buf_2 _287_ (.A(_052_),
    .X(_054_));
 sky130_fd_sc_hd__nor2_1 _288_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .Y(_055_));
 sky130_fd_sc_hd__and3_4 _289_ (.A(_250_),
    .B(_054_),
    .C(_055_),
    .X(_000_));
 sky130_fd_sc_hd__and3_4 _290_ (.A(_253_),
    .B(_054_),
    .C(_055_),
    .X(_007_));
 sky130_fd_sc_hd__and3_4 _291_ (.A(_251_),
    .B(_054_),
    .C(_055_),
    .X(_008_));
 sky130_fd_sc_hd__inv_1 _292_ (.A(_255_),
    .Y(_056_));
 sky130_fd_sc_hd__a211oi_4 _293_ (.A1(_046_),
    .A2(_048_),
    .B1(_051_),
    .C1(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__and2_4 _294_ (.A(_057_),
    .B(_055_),
    .X(_009_));
 sky130_fd_sc_hd__nor2b_1 _295_ (.A(\wr_ptr[3] ),
    .B_N(\wr_ptr[2] ),
    .Y(_058_));
 sky130_fd_sc_hd__and3_4 _296_ (.A(_250_),
    .B(_054_),
    .C(_058_),
    .X(_010_));
 sky130_fd_sc_hd__and3_4 _297_ (.A(_253_),
    .B(_054_),
    .C(_058_),
    .X(_011_));
 sky130_fd_sc_hd__and3_4 _298_ (.A(_251_),
    .B(_054_),
    .C(_058_),
    .X(_012_));
 sky130_fd_sc_hd__and2_4 _299_ (.A(_057_),
    .B(_058_),
    .X(_013_));
 sky130_fd_sc_hd__nor2b_1 _300_ (.A(\wr_ptr[2] ),
    .B_N(\wr_ptr[3] ),
    .Y(_059_));
 sky130_fd_sc_hd__and3_4 _301_ (.A(_250_),
    .B(_054_),
    .C(_059_),
    .X(_014_));
 sky130_fd_sc_hd__and3_4 _302_ (.A(_253_),
    .B(_054_),
    .C(_059_),
    .X(_015_));
 sky130_fd_sc_hd__and3_4 _303_ (.A(_251_),
    .B(_054_),
    .C(_059_),
    .X(_001_));
 sky130_fd_sc_hd__and2_4 _304_ (.A(_057_),
    .B(_059_),
    .X(_002_));
 sky130_fd_sc_hd__inv_1 _305_ (.A(net3),
    .Y(_227_));
 sky130_fd_sc_hd__inv_1 _306_ (.A(_239_),
    .Y(_228_));
 sky130_fd_sc_hd__clkinvlp_4 _307_ (.A(\rd_ptr[3] ),
    .Y(_231_));
 sky130_fd_sc_hd__buf_4 _308_ (.A(\rd_ptr[1] ),
    .X(_060_));
 sky130_fd_sc_hd__inv_2 _309_ (.A(_060_),
    .Y(_224_));
 sky130_fd_sc_hd__inv_1 _310_ (.A(_257_),
    .Y(_225_));
 sky130_fd_sc_hd__buf_4 _311_ (.A(\rd_ptr[2] ),
    .X(_061_));
 sky130_fd_sc_hd__clkinvlp_4 _312_ (.A(_061_),
    .Y(_236_));
 sky130_fd_sc_hd__inv_1 _313_ (.A(\wr_ptr[0] ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_1 _314_ (.A(\wr_ptr[1] ),
    .Y(_249_));
 sky130_fd_sc_hd__clkbuf_4 _315_ (.A(\rd_ptr[0] ),
    .X(_062_));
 sky130_fd_sc_hd__mux4_1 _316_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[4][0] ),
    .A3(\mem[5][0] ),
    .S0(_062_),
    .S1(_061_),
    .X(_063_));
 sky130_fd_sc_hd__nand2_4 _317_ (.A(_231_),
    .B(_224_),
    .Y(_064_));
 sky130_fd_sc_hd__buf_4 _318_ (.A(_060_),
    .X(_065_));
 sky130_fd_sc_hd__nand2_4 _319_ (.A(_231_),
    .B(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__buf_6 _320_ (.A(_062_),
    .X(_067_));
 sky130_fd_sc_hd__buf_6 _321_ (.A(\rd_ptr[2] ),
    .X(_068_));
 sky130_fd_sc_hd__mux4_1 _322_ (.A0(\mem[2][0] ),
    .A1(\mem[3][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_067_),
    .S1(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o22ai_1 _323_ (.A1(_063_),
    .A2(_064_),
    .B1(_066_),
    .B2(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__mux4_1 _324_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S0(_062_),
    .S1(_060_),
    .X(_071_));
 sky130_fd_sc_hd__nand2_8 _325_ (.A(\rd_ptr[3] ),
    .B(_236_),
    .Y(_072_));
 sky130_fd_sc_hd__nand2_8 _326_ (.A(\rd_ptr[3] ),
    .B(_068_),
    .Y(_073_));
 sky130_fd_sc_hd__mux4_1 _327_ (.A0(\mem[12][0] ),
    .A1(\mem[13][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_067_),
    .S1(_065_),
    .X(_074_));
 sky130_fd_sc_hd__o22ai_2 _328_ (.A1(_071_),
    .A2(_072_),
    .B1(_073_),
    .B2(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _329_ (.A(_070_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__o21ai_4 _330_ (.A1(_046_),
    .A2(_049_),
    .B1(net7),
    .Y(_077_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(_076_),
    .A1(net34),
    .S(_077_),
    .X(_019_));
 sky130_fd_sc_hd__buf_4 _332_ (.A(_062_),
    .X(_078_));
 sky130_fd_sc_hd__mux4_1 _333_ (.A0(\mem[2][1] ),
    .A1(\mem[3][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_078_),
    .S1(_061_),
    .X(_079_));
 sky130_fd_sc_hd__buf_6 _334_ (.A(_062_),
    .X(_080_));
 sky130_fd_sc_hd__mux4_1 _335_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[4][1] ),
    .A3(\mem[5][1] ),
    .S0(_080_),
    .S1(_068_),
    .X(_081_));
 sky130_fd_sc_hd__o22ai_1 _336_ (.A1(_066_),
    .A2(_079_),
    .B1(_081_),
    .B2(_064_),
    .Y(_082_));
 sky130_fd_sc_hd__mux4_1 _337_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_080_),
    .S1(_060_),
    .X(_083_));
 sky130_fd_sc_hd__mux4_1 _338_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(_067_),
    .S1(_065_),
    .X(_084_));
 sky130_fd_sc_hd__o22ai_2 _339_ (.A1(_073_),
    .A2(_083_),
    .B1(_084_),
    .B2(_072_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _340_ (.A(_082_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(_086_),
    .A1(net35),
    .S(_077_),
    .X(_020_));
 sky130_fd_sc_hd__mux4_1 _342_ (.A0(\mem[2][2] ),
    .A1(\mem[3][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_078_),
    .S1(_061_),
    .X(_087_));
 sky130_fd_sc_hd__mux4_1 _343_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[4][2] ),
    .A3(\mem[5][2] ),
    .S0(_080_),
    .S1(_068_),
    .X(_088_));
 sky130_fd_sc_hd__o22ai_1 _344_ (.A1(_066_),
    .A2(_087_),
    .B1(_088_),
    .B2(_064_),
    .Y(_089_));
 sky130_fd_sc_hd__mux4_1 _345_ (.A0(\mem[12][2] ),
    .A1(\mem[13][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_080_),
    .S1(_060_),
    .X(_090_));
 sky130_fd_sc_hd__mux4_1 _346_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S0(_067_),
    .S1(_065_),
    .X(_091_));
 sky130_fd_sc_hd__o22ai_1 _347_ (.A1(_073_),
    .A2(_090_),
    .B1(_091_),
    .B2(_072_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _348_ (.A(_089_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(_093_),
    .A1(net36),
    .S(_077_),
    .X(_021_));
 sky130_fd_sc_hd__mux4_1 _350_ (.A0(\mem[2][3] ),
    .A1(\mem[3][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_078_),
    .S1(_061_),
    .X(_094_));
 sky130_fd_sc_hd__mux4_1 _351_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[4][3] ),
    .A3(\mem[5][3] ),
    .S0(_078_),
    .S1(_068_),
    .X(_095_));
 sky130_fd_sc_hd__o22ai_1 _352_ (.A1(_066_),
    .A2(_094_),
    .B1(_095_),
    .B2(_064_),
    .Y(_096_));
 sky130_fd_sc_hd__mux4_2 _353_ (.A0(\mem[12][3] ),
    .A1(\mem[13][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_080_),
    .S1(_060_),
    .X(_097_));
 sky130_fd_sc_hd__mux4_2 _354_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S0(_067_),
    .S1(_065_),
    .X(_098_));
 sky130_fd_sc_hd__o22ai_4 _355_ (.A1(_073_),
    .A2(_097_),
    .B1(_098_),
    .B2(_072_),
    .Y(_099_));
 sky130_fd_sc_hd__nor2_1 _356_ (.A(_096_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(_100_),
    .A1(net37),
    .S(_077_),
    .X(_022_));
 sky130_fd_sc_hd__mux4_1 _358_ (.A0(\mem[2][4] ),
    .A1(\mem[3][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_078_),
    .S1(_061_),
    .X(_101_));
 sky130_fd_sc_hd__mux4_1 _359_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[4][4] ),
    .A3(\mem[5][4] ),
    .S0(_078_),
    .S1(_068_),
    .X(_102_));
 sky130_fd_sc_hd__o22ai_1 _360_ (.A1(_066_),
    .A2(_101_),
    .B1(_102_),
    .B2(_064_),
    .Y(_103_));
 sky130_fd_sc_hd__mux4_1 _361_ (.A0(\mem[12][4] ),
    .A1(\mem[13][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_080_),
    .S1(_060_),
    .X(_104_));
 sky130_fd_sc_hd__mux4_1 _362_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[11][4] ),
    .S0(_067_),
    .S1(_065_),
    .X(_105_));
 sky130_fd_sc_hd__o22ai_2 _363_ (.A1(_073_),
    .A2(_104_),
    .B1(_105_),
    .B2(_072_),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _364_ (.A(_103_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(_107_),
    .A1(net38),
    .S(_077_),
    .X(_023_));
 sky130_fd_sc_hd__mux4_1 _366_ (.A0(\mem[2][5] ),
    .A1(\mem[3][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_078_),
    .S1(_061_),
    .X(_108_));
 sky130_fd_sc_hd__mux4_1 _367_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[4][5] ),
    .A3(\mem[5][5] ),
    .S0(_078_),
    .S1(_068_),
    .X(_109_));
 sky130_fd_sc_hd__o22ai_1 _368_ (.A1(_066_),
    .A2(_108_),
    .B1(_109_),
    .B2(_064_),
    .Y(_110_));
 sky130_fd_sc_hd__mux4_2 _369_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_080_),
    .S1(_060_),
    .X(_111_));
 sky130_fd_sc_hd__mux4_2 _370_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(_067_),
    .S1(_065_),
    .X(_112_));
 sky130_fd_sc_hd__o22ai_4 _371_ (.A1(_073_),
    .A2(_111_),
    .B1(_112_),
    .B2(_072_),
    .Y(_113_));
 sky130_fd_sc_hd__nor2_1 _372_ (.A(_110_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(_114_),
    .A1(net39),
    .S(_077_),
    .X(_024_));
 sky130_fd_sc_hd__mux4_1 _374_ (.A0(\mem[2][6] ),
    .A1(\mem[3][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_062_),
    .S1(_061_),
    .X(_115_));
 sky130_fd_sc_hd__mux4_1 _375_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[4][6] ),
    .A3(\mem[5][6] ),
    .S0(_078_),
    .S1(_068_),
    .X(_116_));
 sky130_fd_sc_hd__o22ai_1 _376_ (.A1(_066_),
    .A2(_115_),
    .B1(_116_),
    .B2(_064_),
    .Y(_117_));
 sky130_fd_sc_hd__mux4_1 _377_ (.A0(\mem[12][6] ),
    .A1(\mem[13][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_080_),
    .S1(_060_),
    .X(_118_));
 sky130_fd_sc_hd__mux4_1 _378_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[10][6] ),
    .A3(\mem[11][6] ),
    .S0(_067_),
    .S1(_065_),
    .X(_119_));
 sky130_fd_sc_hd__o22ai_4 _379_ (.A1(_073_),
    .A2(_118_),
    .B1(_119_),
    .B2(_072_),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_1 _380_ (.A(_117_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(_121_),
    .A1(net40),
    .S(_077_),
    .X(_025_));
 sky130_fd_sc_hd__mux4_1 _382_ (.A0(\mem[2][7] ),
    .A1(\mem[3][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_062_),
    .S1(_061_),
    .X(_122_));
 sky130_fd_sc_hd__mux4_1 _383_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[4][7] ),
    .A3(\mem[5][7] ),
    .S0(_078_),
    .S1(_061_),
    .X(_123_));
 sky130_fd_sc_hd__o22ai_1 _384_ (.A1(_066_),
    .A2(_122_),
    .B1(_123_),
    .B2(_064_),
    .Y(_124_));
 sky130_fd_sc_hd__mux4_1 _385_ (.A0(\mem[12][7] ),
    .A1(\mem[13][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_080_),
    .S1(_060_),
    .X(_125_));
 sky130_fd_sc_hd__mux4_1 _386_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[10][7] ),
    .A3(\mem[11][7] ),
    .S0(_080_),
    .S1(_065_),
    .X(_126_));
 sky130_fd_sc_hd__o22ai_2 _387_ (.A1(_073_),
    .A2(_125_),
    .B1(_126_),
    .B2(_072_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _388_ (.A(_124_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(_128_),
    .A1(net41),
    .S(_077_),
    .X(_026_));
 sky130_fd_sc_hd__xnor2_1 _390_ (.A(_067_),
    .B(_077_),
    .Y(_027_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(_018_),
    .A1(_065_),
    .S(_077_),
    .X(_028_));
 sky130_fd_sc_hd__o211ai_1 _392_ (.A1(net24),
    .A2(_049_),
    .B1(net7),
    .C1(_248_),
    .Y(_129_));
 sky130_fd_sc_hd__xnor2_1 _393_ (.A(_068_),
    .B(_129_),
    .Y(_029_));
 sky130_fd_sc_hd__nand2_1 _394_ (.A(net7),
    .B(_067_),
    .Y(_130_));
 sky130_fd_sc_hd__nor3_1 _395_ (.A(_224_),
    .B(_236_),
    .C(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__o21ai_0 _396_ (.A1(net24),
    .A2(_049_),
    .B1(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__xnor2_1 _397_ (.A(\rd_ptr[3] ),
    .B(_132_),
    .Y(_030_));
 sky130_fd_sc_hd__and4_1 _398_ (.A(net7),
    .B(\rd_ptr[3] ),
    .C(_068_),
    .D(_248_),
    .X(_133_));
 sky130_fd_sc_hd__o21ai_1 _399_ (.A1(net24),
    .A2(_049_),
    .B1(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__xnor2_1 _400_ (.A(\rd_ptr[4] ),
    .B(_134_),
    .Y(_031_));
 sky130_fd_sc_hd__xnor2_1 _401_ (.A(_016_),
    .B(_054_),
    .Y(_032_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\wr_ptr[1] ),
    .A1(_017_),
    .S(_052_),
    .X(_033_));
 sky130_fd_sc_hd__xor2_1 _403_ (.A(\wr_ptr[2] ),
    .B(_057_),
    .X(_034_));
 sky130_fd_sc_hd__nand4_1 _404_ (.A(net16),
    .B(\wr_ptr[2] ),
    .C(\wr_ptr[1] ),
    .D(\wr_ptr[0] ),
    .Y(_135_));
 sky130_fd_sc_hd__a21oi_1 _405_ (.A1(net24),
    .A2(_048_),
    .B1(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__xor2_1 _406_ (.A(\wr_ptr[3] ),
    .B(_136_),
    .X(_035_));
 sky130_fd_sc_hd__xor2_1 _407_ (.A(\wr_ptr[4] ),
    .B(_006_),
    .X(_036_));
 sky130_fd_sc_hd__xor2_1 _408_ (.A(_258_),
    .B(net21),
    .X(_137_));
 sky130_fd_sc_hd__nor4_1 _409_ (.A(net23),
    .B(net22),
    .C(net24),
    .D(_137_),
    .Y(net17));
 sky130_fd_sc_hd__nand3_1 _410_ (.A(net21),
    .B(net23),
    .C(net22),
    .Y(_138_));
 sky130_fd_sc_hd__nand2_1 _411_ (.A(net24),
    .B(_049_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_0 _412_ (.A1(net24),
    .A2(_138_),
    .B1(_139_),
    .Y(net18));
 sky130_fd_sc_hd__a21o_1 _413_ (.A1(_239_),
    .A2(_242_),
    .B1(_241_),
    .X(_140_));
 sky130_fd_sc_hd__a21oi_2 _414_ (.A1(_244_),
    .A2(_140_),
    .B1(_243_),
    .Y(_141_));
 sky130_fd_sc_hd__xnor2_2 _415_ (.A(net5),
    .B(\rd_ptr[3] ),
    .Y(_142_));
 sky130_fd_sc_hd__xnor2_4 _416_ (.A(_141_),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__clkbuf_4 _417_ (.A(_143_),
    .X(_144_));
 sky130_fd_sc_hd__buf_2 _418_ (.A(_240_),
    .X(_145_));
 sky130_fd_sc_hd__buf_6 _419_ (.A(_145_),
    .X(_146_));
 sky130_fd_sc_hd__clkbuf_8 _420_ (.A(_146_),
    .X(_147_));
 sky130_fd_sc_hd__buf_4 _421_ (.A(_230_),
    .X(_148_));
 sky130_fd_sc_hd__buf_4 _422_ (.A(_148_),
    .X(_149_));
 sky130_fd_sc_hd__mux4_1 _423_ (.A0(\mem[4][0] ),
    .A1(\mem[5][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_147_),
    .S1(_149_),
    .X(_150_));
 sky130_fd_sc_hd__mux4_1 _424_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[2][0] ),
    .A3(\mem[3][0] ),
    .S0(_147_),
    .S1(_149_),
    .X(_151_));
 sky130_fd_sc_hd__xor2_4 _425_ (.A(_229_),
    .B(_244_),
    .X(_152_));
 sky130_fd_sc_hd__buf_8 _426_ (.A(_152_),
    .X(_153_));
 sky130_fd_sc_hd__buf_6 _427_ (.A(_153_),
    .X(_154_));
 sky130_fd_sc_hd__mux2i_2 _428_ (.A0(_150_),
    .A1(_151_),
    .S(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__buf_6 _429_ (.A(_145_),
    .X(_156_));
 sky130_fd_sc_hd__buf_6 _430_ (.A(_230_),
    .X(_157_));
 sky130_fd_sc_hd__mux4_1 _431_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S0(_156_),
    .S1(_157_),
    .X(_158_));
 sky130_fd_sc_hd__mux4_1 _432_ (.A0(\mem[12][0] ),
    .A1(\mem[13][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_146_),
    .S1(_148_),
    .X(_159_));
 sky130_fd_sc_hd__nor2b_1 _433_ (.A(_153_),
    .B_N(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__a211oi_1 _434_ (.A1(_154_),
    .A2(_158_),
    .B1(_160_),
    .C1(_144_),
    .Y(_161_));
 sky130_fd_sc_hd__nand2_1 _435_ (.A(_037_),
    .B(_038_),
    .Y(_162_));
 sky130_fd_sc_hd__and2_0 _436_ (.A(_233_),
    .B(net5),
    .X(_163_));
 sky130_fd_sc_hd__nor3_1 _437_ (.A(_258_),
    .B(_246_),
    .C(net2),
    .Y(_164_));
 sky130_fd_sc_hd__o21ai_0 _438_ (.A1(_246_),
    .A2(_247_),
    .B1(net4),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_0 _439_ (.A1(_164_),
    .A2(_165_),
    .B1(net22),
    .Y(_166_));
 sky130_fd_sc_hd__o21ai_0 _440_ (.A1(_258_),
    .A2(net2),
    .B1(_247_),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(net4),
    .B(_246_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _442_ (.A(_167_),
    .B(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__nor4b_1 _443_ (.A(_233_),
    .B(_040_),
    .C(_041_),
    .D_N(net5),
    .Y(_170_));
 sky130_fd_sc_hd__a221oi_2 _444_ (.A1(_162_),
    .A2(_163_),
    .B1(_166_),
    .B2(_169_),
    .C1(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__a211oi_2 _445_ (.A1(_037_),
    .A2(_038_),
    .B1(_233_),
    .C1(net5),
    .Y(_172_));
 sky130_fd_sc_hd__nor3b_1 _446_ (.A(net5),
    .B(_162_),
    .C_N(_233_),
    .Y(_173_));
 sky130_fd_sc_hd__o41ai_4 _447_ (.A1(_046_),
    .A2(_171_),
    .A3(_172_),
    .A4(_173_),
    .B1(net6),
    .Y(_174_));
 sky130_fd_sc_hd__a211oi_1 _448_ (.A1(_144_),
    .A2(_155_),
    .B1(_161_),
    .C1(_174_),
    .Y(net26));
 sky130_fd_sc_hd__mux4_1 _449_ (.A0(\mem[4][1] ),
    .A1(\mem[5][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_147_),
    .S1(_149_),
    .X(_175_));
 sky130_fd_sc_hd__mux4_1 _450_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[2][1] ),
    .A3(\mem[3][1] ),
    .S0(_147_),
    .S1(_149_),
    .X(_176_));
 sky130_fd_sc_hd__mux2i_2 _451_ (.A0(_175_),
    .A1(_176_),
    .S(_154_),
    .Y(_177_));
 sky130_fd_sc_hd__mux4_1 _452_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(_156_),
    .S1(_157_),
    .X(_178_));
 sky130_fd_sc_hd__mux4_1 _453_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_146_),
    .S1(_148_),
    .X(_179_));
 sky130_fd_sc_hd__nor2b_1 _454_ (.A(_153_),
    .B_N(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__a211oi_1 _455_ (.A1(_154_),
    .A2(_178_),
    .B1(_180_),
    .C1(_144_),
    .Y(_181_));
 sky130_fd_sc_hd__a211oi_1 _456_ (.A1(_144_),
    .A2(_177_),
    .B1(_181_),
    .C1(_174_),
    .Y(net27));
 sky130_fd_sc_hd__mux4_1 _457_ (.A0(\mem[4][2] ),
    .A1(\mem[5][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_147_),
    .S1(_149_),
    .X(_182_));
 sky130_fd_sc_hd__mux4_1 _458_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[2][2] ),
    .A3(\mem[3][2] ),
    .S0(_156_),
    .S1(_157_),
    .X(_183_));
 sky130_fd_sc_hd__mux2i_1 _459_ (.A0(_182_),
    .A1(_183_),
    .S(_153_),
    .Y(_184_));
 sky130_fd_sc_hd__mux4_1 _460_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S0(_156_),
    .S1(_157_),
    .X(_185_));
 sky130_fd_sc_hd__mux4_1 _461_ (.A0(\mem[12][2] ),
    .A1(\mem[13][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_146_),
    .S1(_148_),
    .X(_186_));
 sky130_fd_sc_hd__nor2b_1 _462_ (.A(_153_),
    .B_N(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a211oi_1 _463_ (.A1(_154_),
    .A2(_185_),
    .B1(_187_),
    .C1(_143_),
    .Y(_188_));
 sky130_fd_sc_hd__a211oi_2 _464_ (.A1(_144_),
    .A2(_184_),
    .B1(_188_),
    .C1(_174_),
    .Y(net28));
 sky130_fd_sc_hd__mux4_1 _465_ (.A0(\mem[4][3] ),
    .A1(\mem[5][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_147_),
    .S1(_149_),
    .X(_189_));
 sky130_fd_sc_hd__mux4_1 _466_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[2][3] ),
    .A3(\mem[3][3] ),
    .S0(_156_),
    .S1(_157_),
    .X(_190_));
 sky130_fd_sc_hd__mux2i_4 _467_ (.A0(_189_),
    .A1(_190_),
    .S(_153_),
    .Y(_191_));
 sky130_fd_sc_hd__mux4_1 _468_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S0(_156_),
    .S1(_157_),
    .X(_192_));
 sky130_fd_sc_hd__mux4_1 _469_ (.A0(\mem[12][3] ),
    .A1(\mem[13][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_146_),
    .S1(_148_),
    .X(_193_));
 sky130_fd_sc_hd__nor2b_1 _470_ (.A(_152_),
    .B_N(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__a211oi_1 _471_ (.A1(_154_),
    .A2(_192_),
    .B1(_194_),
    .C1(_143_),
    .Y(_195_));
 sky130_fd_sc_hd__a211oi_2 _472_ (.A1(_144_),
    .A2(_191_),
    .B1(_195_),
    .C1(_174_),
    .Y(net29));
 sky130_fd_sc_hd__mux4_1 _473_ (.A0(\mem[4][4] ),
    .A1(\mem[5][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_147_),
    .S1(_149_),
    .X(_196_));
 sky130_fd_sc_hd__mux4_1 _474_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[2][4] ),
    .A3(\mem[3][4] ),
    .S0(_156_),
    .S1(_157_),
    .X(_197_));
 sky130_fd_sc_hd__mux2i_2 _475_ (.A0(_196_),
    .A1(_197_),
    .S(_153_),
    .Y(_198_));
 sky130_fd_sc_hd__mux4_1 _476_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[11][4] ),
    .S0(_146_),
    .S1(_148_),
    .X(_199_));
 sky130_fd_sc_hd__mux4_1 _477_ (.A0(\mem[12][4] ),
    .A1(\mem[13][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_146_),
    .S1(_148_),
    .X(_200_));
 sky130_fd_sc_hd__nor2b_1 _478_ (.A(_152_),
    .B_N(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__a211oi_2 _479_ (.A1(_154_),
    .A2(_199_),
    .B1(_201_),
    .C1(_143_),
    .Y(_202_));
 sky130_fd_sc_hd__a211oi_2 _480_ (.A1(_144_),
    .A2(_198_),
    .B1(_202_),
    .C1(_174_),
    .Y(net30));
 sky130_fd_sc_hd__mux4_1 _481_ (.A0(\mem[4][5] ),
    .A1(\mem[5][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_147_),
    .S1(_149_),
    .X(_203_));
 sky130_fd_sc_hd__mux4_1 _482_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[2][5] ),
    .A3(\mem[3][5] ),
    .S0(_156_),
    .S1(_157_),
    .X(_204_));
 sky130_fd_sc_hd__mux2i_4 _483_ (.A0(_203_),
    .A1(_204_),
    .S(_153_),
    .Y(_205_));
 sky130_fd_sc_hd__mux4_1 _484_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(_146_),
    .S1(_148_),
    .X(_206_));
 sky130_fd_sc_hd__mux4_1 _485_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_145_),
    .S1(_230_),
    .X(_207_));
 sky130_fd_sc_hd__nor2b_1 _486_ (.A(_152_),
    .B_N(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__a211oi_1 _487_ (.A1(_154_),
    .A2(_206_),
    .B1(_208_),
    .C1(_143_),
    .Y(_209_));
 sky130_fd_sc_hd__a211oi_1 _488_ (.A1(_144_),
    .A2(_205_),
    .B1(_209_),
    .C1(_174_),
    .Y(net31));
 sky130_fd_sc_hd__mux4_1 _489_ (.A0(\mem[4][6] ),
    .A1(\mem[5][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_147_),
    .S1(_149_),
    .X(_210_));
 sky130_fd_sc_hd__mux4_1 _490_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[2][6] ),
    .A3(\mem[3][6] ),
    .S0(_156_),
    .S1(_157_),
    .X(_211_));
 sky130_fd_sc_hd__mux2i_2 _491_ (.A0(_210_),
    .A1(_211_),
    .S(_153_),
    .Y(_212_));
 sky130_fd_sc_hd__mux4_1 _492_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[10][6] ),
    .A3(\mem[11][6] ),
    .S0(_146_),
    .S1(_148_),
    .X(_213_));
 sky130_fd_sc_hd__mux4_1 _493_ (.A0(\mem[12][6] ),
    .A1(\mem[13][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_145_),
    .S1(_230_),
    .X(_214_));
 sky130_fd_sc_hd__nor2b_1 _494_ (.A(_152_),
    .B_N(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__a211oi_1 _495_ (.A1(_154_),
    .A2(_213_),
    .B1(_215_),
    .C1(_143_),
    .Y(_216_));
 sky130_fd_sc_hd__a211oi_1 _496_ (.A1(_144_),
    .A2(_212_),
    .B1(_216_),
    .C1(_174_),
    .Y(net32));
 sky130_fd_sc_hd__mux4_1 _497_ (.A0(\mem[4][7] ),
    .A1(\mem[5][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_147_),
    .S1(_149_),
    .X(_217_));
 sky130_fd_sc_hd__mux4_1 _498_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[2][7] ),
    .A3(\mem[3][7] ),
    .S0(_156_),
    .S1(_157_),
    .X(_218_));
 sky130_fd_sc_hd__mux2i_2 _499_ (.A0(_217_),
    .A1(_218_),
    .S(_153_),
    .Y(_219_));
 sky130_fd_sc_hd__mux4_1 _500_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[10][7] ),
    .A3(\mem[11][7] ),
    .S0(_146_),
    .S1(_148_),
    .X(_220_));
 sky130_fd_sc_hd__mux4_1 _501_ (.A0(\mem[12][7] ),
    .A1(\mem[13][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_145_),
    .S1(_230_),
    .X(_221_));
 sky130_fd_sc_hd__nor2b_1 _502_ (.A(_152_),
    .B_N(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__a211oi_1 _503_ (.A1(_154_),
    .A2(_220_),
    .B1(_222_),
    .C1(_143_),
    .Y(_223_));
 sky130_fd_sc_hd__a211oi_1 _504_ (.A1(_144_),
    .A2(_219_),
    .B1(_223_),
    .C1(_174_),
    .Y(net33));
 sky130_fd_sc_hd__fa_2 _505_ (.A(_224_),
    .B(\wr_ptr[1] ),
    .CIN(_225_),
    .COUT(_226_),
    .SUM(net21));
 sky130_fd_sc_hd__fa_4 _506_ (.A(_227_),
    .B(_224_),
    .CIN(_228_),
    .COUT(_229_),
    .SUM(_230_));
 sky130_fd_sc_hd__ha_2 _507_ (.A(_231_),
    .B(\wr_ptr[3] ),
    .COUT(_232_),
    .SUM(_233_));
 sky130_fd_sc_hd__ha_1 _508_ (.A(_224_),
    .B(\wr_ptr[1] ),
    .COUT(_234_),
    .SUM(_235_));
 sky130_fd_sc_hd__ha_2 _509_ (.A(_236_),
    .B(\wr_ptr[2] ),
    .COUT(_237_),
    .SUM(_238_));
 sky130_fd_sc_hd__ha_1 _510_ (.A(net2),
    .B(\rd_ptr[0] ),
    .COUT(_239_),
    .SUM(_240_));
 sky130_fd_sc_hd__ha_1 _511_ (.A(net3),
    .B(\rd_ptr[1] ),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__ha_2 _512_ (.A(net4),
    .B(\rd_ptr[2] ),
    .COUT(_243_),
    .SUM(_244_));
 sky130_fd_sc_hd__ha_1 _513_ (.A(net3),
    .B(_245_),
    .COUT(_246_),
    .SUM(_247_));
 sky130_fd_sc_hd__ha_1 _514_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_248_),
    .SUM(_018_));
 sky130_fd_sc_hd__ha_1 _515_ (.A(_016_),
    .B(_249_),
    .COUT(_250_),
    .SUM(_017_));
 sky130_fd_sc_hd__ha_1 _516_ (.A(_016_),
    .B(\wr_ptr[1] ),
    .COUT(_251_),
    .SUM(_252_));
 sky130_fd_sc_hd__ha_1 _517_ (.A(\wr_ptr[0] ),
    .B(_249_),
    .COUT(_253_),
    .SUM(_254_));
 sky130_fd_sc_hd__ha_1 _518_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__ha_1 _519_ (.A(\rd_ptr[0] ),
    .B(_016_),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net10),
    .DE(_000_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net11),
    .DE(_000_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net12),
    .DE(_000_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net13),
    .DE(_000_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net14),
    .DE(_000_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net15),
    .DE(_000_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net11),
    .DE(_001_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net12),
    .DE(_001_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net13),
    .DE(_001_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net14),
    .DE(_001_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net15),
    .DE(_001_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net11),
    .DE(_002_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net12),
    .DE(_002_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net13),
    .DE(_002_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net14),
    .DE(_002_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net15),
    .DE(_002_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net11),
    .DE(_003_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net12),
    .DE(_003_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net13),
    .DE(_003_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net14),
    .DE(_003_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net15),
    .DE(_003_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net11),
    .DE(_004_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net12),
    .DE(_004_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net13),
    .DE(_004_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net14),
    .DE(_004_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net15),
    .DE(_004_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net11),
    .DE(_005_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net12),
    .DE(_005_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net13),
    .DE(_005_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net14),
    .DE(_005_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net15),
    .DE(_005_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net11),
    .DE(_006_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net12),
    .DE(_006_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net13),
    .DE(_006_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net14),
    .DE(_006_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net15),
    .DE(_006_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net11),
    .DE(_007_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net12),
    .DE(_007_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net13),
    .DE(_007_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net14),
    .DE(_007_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net15),
    .DE(_007_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net11),
    .DE(_008_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net12),
    .DE(_008_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net13),
    .DE(_008_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net14),
    .DE(_008_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net15),
    .DE(_008_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net11),
    .DE(_009_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net12),
    .DE(_009_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net13),
    .DE(_009_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net14),
    .DE(_009_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net15),
    .DE(_009_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net11),
    .DE(_010_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net12),
    .DE(_010_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net13),
    .DE(_010_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net14),
    .DE(_010_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net15),
    .DE(_010_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net12),
    .DE(_011_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net13),
    .DE(_011_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net14),
    .DE(_011_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net15),
    .DE(_011_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net12),
    .DE(_012_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net13),
    .DE(_012_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net14),
    .DE(_012_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net15),
    .DE(_012_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net12),
    .DE(_013_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net13),
    .DE(_013_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net14),
    .DE(_013_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net15),
    .DE(_013_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net12),
    .DE(_014_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net13),
    .DE(_014_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net14),
    .DE(_014_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net15),
    .DE(_014_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net12),
    .DE(_015_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net13),
    .DE(_015_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net14),
    .DE(_015_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net15),
    .DE(_015_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[0]$_DFFE_PN0P_  (.D(_019_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[1]$_DFFE_PN0P_  (.D(_020_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[2]$_DFFE_PN0P_  (.D(_021_),
    .Q(net36),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[3]$_DFFE_PN0P_  (.D(_022_),
    .Q(net37),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[4]$_DFFE_PN0P_  (.D(_023_),
    .Q(net38),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[5]$_DFFE_PN0P_  (.D(_024_),
    .Q(net39),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[6]$_DFFE_PN0P_  (.D(_025_),
    .Q(net40),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[7]$_DFFE_PN0P_  (.D(_026_),
    .Q(net41),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_027_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_028_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_029_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr[3]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_032_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_033_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[2]$_DFFE_PN0P_  (.D(_034_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[3]$_DFFE_PN0P_  (.D(_035_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_036_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__buf_8 hold1 (.A(net42),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_224 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(peek_addr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(peek_addr[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(peek_addr[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(peek_addr[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(peek_en),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(rd_en),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[0]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(wr_data[1]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input10 (.A(wr_data[3]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input11 (.A(wr_data[4]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input12 (.A(wr_data[5]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input13 (.A(wr_data[6]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input14 (.A(wr_data[7]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(wr_en),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(fifo_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(fifo_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(fifo_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(fifo_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(fifo_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(peek_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(peek_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(peek_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(peek_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(peek_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(peek_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(peek_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(peek_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net42));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_289 ();
endmodule
