module pwm_generator (clk,
    enable,
    pwm_out,
    rst_n,
    duty_cycle,
    period);
 input clk;
 input enable;
 output pwm_out;
 input rst_n;
 input [7:0] duty_cycle;
 input [7:0] period;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \duty_reg[0] ;
 wire \duty_reg[1] ;
 wire \duty_reg[2] ;
 wire \duty_reg[3] ;
 wire \duty_reg[4] ;
 wire \duty_reg[5] ;
 wire \duty_reg[6] ;
 wire \duty_reg[7] ;
 wire \period_reg[0] ;
 wire \period_reg[1] ;
 wire \period_reg[2] ;
 wire \period_reg[3] ;
 wire \period_reg[4] ;
 wire \period_reg[5] ;
 wire \period_reg[6] ;
 wire \period_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _117_ (.I(\counter[1] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _118_ (.I(\counter[3] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _119_ (.I(\counter[2] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _120_ (.I(\counter[7] ),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _121_ (.I(\counter[6] ),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _122_ (.I(\counter[5] ),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _123_ (.I(\counter[4] ),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _124_ (.I(\period_reg[0] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _125_ (.I(\duty_reg[7] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _126_ (.I(\duty_reg[6] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _127_ (.I(\duty_reg[5] ),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _128_ (.I(\duty_reg[4] ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _129_ (.I(\duty_reg[3] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _130_ (.I(\duty_reg[2] ),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _131_ (.I(\duty_reg[1] ),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _132_ (.I(net10),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _133_ (.I(_025_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _134_ (.A1(_078_),
    .A2(_081_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_071_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _136_ (.A1(_075_),
    .A2(_028_),
    .B(_074_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _137_ (.A1(_078_),
    .A2(_080_),
    .B(_077_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _138_ (.A1(_027_),
    .A2(_029_),
    .B(_030_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _139_ (.A1(_084_),
    .A2(_093_),
    .A3(_090_),
    .A4(_087_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _140_ (.A1(_075_),
    .A2(_078_),
    .A3(_072_),
    .A4(_081_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _141_ (.A1(_032_),
    .A2(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _142_ (.A1(_032_),
    .A2(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _143_ (.A1(_090_),
    .A2(_092_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _144_ (.A1(_089_),
    .A2(_036_),
    .B(_084_),
    .C(_087_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _145_ (.A1(_084_),
    .A2(_086_),
    .B(_083_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _146_ (.A1(_032_),
    .A2(_033_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _147_ (.A1(_037_),
    .A2(_038_),
    .B(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _148_ (.A1(_031_),
    .A2(_035_),
    .B(_040_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _149_ (.A1(_026_),
    .A2(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _150_ (.I(\counter[0] ),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(_026_),
    .I1(_042_),
    .S(_043_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _152_ (.A1(_095_),
    .A2(_025_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _153_ (.A1(_073_),
    .A2(_025_),
    .B1(_041_),
    .B2(_044_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _154_ (.A1(_094_),
    .A2(_079_),
    .A3(_025_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _155_ (.A1(_094_),
    .A2(_079_),
    .A3(_041_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _156_ (.A1(_079_),
    .A2(_025_),
    .B1(_041_),
    .B2(_045_),
    .C(_046_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _157_ (.A1(_076_),
    .A2(_025_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _158_ (.A1(\counter[0] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(_076_),
    .I1(_047_),
    .S(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _160_ (.A1(_076_),
    .A2(_025_),
    .B1(_041_),
    .B2(_049_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _161_ (.A1(_025_),
    .A2(_041_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _162_ (.A1(_094_),
    .A2(\counter[2] ),
    .A3(\counter[3] ),
    .A4(net10),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _163_ (.A1(_091_),
    .A2(_051_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _164_ (.A1(_050_),
    .A2(_052_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _165_ (.A1(\counter[3] ),
    .A2(\counter[4] ),
    .A3(_025_),
    .A4(_048_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _166_ (.A1(_088_),
    .A2(_053_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _167_ (.A1(_050_),
    .A2(_054_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _168_ (.A1(\counter[4] ),
    .A2(\counter[5] ),
    .A3(_051_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _169_ (.A1(_085_),
    .A2(_055_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _170_ (.A1(_050_),
    .A2(_056_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _171_ (.A1(\counter[5] ),
    .A2(\counter[6] ),
    .A3(_053_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _172_ (.A1(_082_),
    .A2(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _173_ (.A1(_050_),
    .A2(_058_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _174_ (.I(_039_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _175_ (.I0(\duty_reg[0] ),
    .I1(net2),
    .S(_059_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _176_ (.I0(\duty_reg[1] ),
    .I1(net3),
    .S(_059_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _177_ (.I0(\duty_reg[2] ),
    .I1(net4),
    .S(_059_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _178_ (.I0(\duty_reg[3] ),
    .I1(net5),
    .S(_059_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _179_ (.I0(\duty_reg[4] ),
    .I1(net6),
    .S(_059_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _180_ (.I0(\duty_reg[5] ),
    .I1(net7),
    .S(_059_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _181_ (.I0(\duty_reg[6] ),
    .I1(net8),
    .S(_059_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _182_ (.I0(\duty_reg[7] ),
    .I1(net9),
    .S(_059_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _183_ (.I0(\period_reg[0] ),
    .I1(net11),
    .S(_059_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _184_ (.I0(\period_reg[1] ),
    .I1(net12),
    .S(_059_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _185_ (.I0(\period_reg[2] ),
    .I1(net13),
    .S(_039_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _186_ (.I0(\period_reg[3] ),
    .I1(net14),
    .S(_039_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _187_ (.I0(\period_reg[4] ),
    .I1(net15),
    .S(_039_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _188_ (.I0(\period_reg[5] ),
    .I1(net16),
    .S(_039_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _189_ (.I0(\period_reg[6] ),
    .I1(net17),
    .S(_039_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _190_ (.I0(\period_reg[7] ),
    .I1(net18),
    .S(_039_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _191_ (.I(_103_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _192_ (.A1(_106_),
    .A2(_107_),
    .B(_104_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _193_ (.A1(_060_),
    .A2(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _194_ (.A1(_098_),
    .A2(_101_),
    .A3(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _195_ (.A1(_043_),
    .A2(\duty_reg[0] ),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _196_ (.A1(_116_),
    .A2(_064_),
    .B(_115_),
    .C(_112_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _197_ (.A1(_113_),
    .A2(_112_),
    .B(_110_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _198_ (.A1(_106_),
    .A2(_104_),
    .B(_103_),
    .C(_109_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _199_ (.A1(_065_),
    .A2(_066_),
    .B(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _200_ (.A1(_098_),
    .A2(_100_),
    .B1(_063_),
    .B2(_068_),
    .C(_097_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _201_ (.I0(net20),
    .I1(_069_),
    .S(_025_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _202_ (.A(\counter[0] ),
    .B(_070_),
    .CO(_071_),
    .S(_072_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _203_ (.A(_073_),
    .B(\period_reg[1] ),
    .CO(_074_),
    .S(_075_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _204_ (.A(_076_),
    .B(\period_reg[3] ),
    .CO(_077_),
    .S(_078_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _205_ (.A(_079_),
    .B(\period_reg[2] ),
    .CO(_080_),
    .S(_081_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _206_ (.A(_082_),
    .B(\period_reg[7] ),
    .CO(_083_),
    .S(_084_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _207_ (.A(_085_),
    .B(\period_reg[6] ),
    .CO(_086_),
    .S(_087_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _208_ (.A(_088_),
    .B(\period_reg[5] ),
    .CO(_089_),
    .S(_090_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _209_ (.A(_091_),
    .B(\period_reg[4] ),
    .CO(_092_),
    .S(_093_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _210_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_094_),
    .S(_095_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _211_ (.A(\counter[7] ),
    .B(_096_),
    .CO(_097_),
    .S(_098_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _212_ (.A(\counter[6] ),
    .B(_099_),
    .CO(_100_),
    .S(_101_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _213_ (.A(\counter[5] ),
    .B(_102_),
    .CO(_103_),
    .S(_104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _214_ (.A(\counter[4] ),
    .B(_105_),
    .CO(_106_),
    .S(_107_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _215_ (.A(\counter[3] ),
    .B(_108_),
    .CO(_109_),
    .S(_110_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _216_ (.A(\counter[2] ),
    .B(_111_),
    .CO(_112_),
    .S(_113_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _217_ (.A(\counter[1] ),
    .B(_114_),
    .CO(_115_),
    .S(_116_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[3]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[4]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[5]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[6]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter[7]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[0]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[1]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[2]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[3]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[4]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[5]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \duty_reg[6]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \duty_reg[7]$_DFFE_PN1P_  (.D(_015_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\duty_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[0]$_DFFE_PN1P_  (.D(_016_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[1]$_DFFE_PN1P_  (.D(_017_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[2]$_DFFE_PN1P_  (.D(_018_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[3]$_DFFE_PN1P_  (.D(_019_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[4]$_DFFE_PN1P_  (.D(_020_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[5]$_DFFE_PN1P_  (.D(_021_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[6]$_DFFE_PN1P_  (.D(_022_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \period_reg[7]$_DFFE_PN1P_  (.D(_023_),
    .SETN(net19),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\period_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \pwm_out$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 hold1 (.I(net19),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_145 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(duty_cycle[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(duty_cycle[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(duty_cycle[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(duty_cycle[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(duty_cycle[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(duty_cycle[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(duty_cycle[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(duty_cycle[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(enable),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(period[0]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(period[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(period[2]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(period[3]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(period[4]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(period[5]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(period[6]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(period[7]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input18 (.I(rst_n),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(pwm_out));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_442 ();
endmodule
