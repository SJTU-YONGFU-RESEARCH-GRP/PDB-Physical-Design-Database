module non_restoring_divider (busy,
    clk,
    error,
    rst_n,
    start,
    valid,
    dividend,
    divisor,
    quotient,
    remainder);
 output busy;
 input clk;
 output error;
 input rst_n;
 input start;
 output valid;
 input [7:0] dividend;
 input [7:0] divisor;
 output [7:0] quotient;
 output [7:0] remainder;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire \div_reg[0] ;
 wire \div_reg[1] ;
 wire \div_reg[2] ;
 wire \div_reg[3] ;
 wire \div_reg[4] ;
 wire \div_reg[5] ;
 wire \div_reg[6] ;
 wire \div_reg[7] ;
 wire \iter[0] ;
 wire \iter[1] ;
 wire \iter[2] ;
 wire \iter[3] ;
 wire \quot[0] ;
 wire \quot[1] ;
 wire \quot[2] ;
 wire \quot[3] ;
 wire \quot[4] ;
 wire \quot[5] ;
 wire \quot[6] ;
 wire \quot[7] ;
 wire \rem[0] ;
 wire \rem[1] ;
 wire \rem[2] ;
 wire \rem[3] ;
 wire \rem[4] ;
 wire \rem[5] ;
 wire \rem[6] ;
 wire \rem[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X1 _339_ (.A(rst_n),
    .Z(_051_));
 INV_X2 _340_ (.A(_051_),
    .ZN(_052_));
 CLKBUF_X3 _341_ (.A(_052_),
    .Z(_053_));
 CLKBUF_X3 _342_ (.A(\state[0] ),
    .Z(_054_));
 CLKBUF_X2 _343_ (.A(start),
    .Z(_055_));
 INV_X1 _344_ (.A(_055_),
    .ZN(_056_));
 NOR4_X4 _345_ (.A1(net14),
    .A2(net13),
    .A3(net16),
    .A4(net15),
    .ZN(_057_));
 NOR4_X4 _346_ (.A1(net10),
    .A2(net9),
    .A3(net12),
    .A4(net11),
    .ZN(_058_));
 AOI21_X4 _347_ (.A(_056_),
    .B1(_057_),
    .B2(_058_),
    .ZN(_059_));
 NAND2_X1 _348_ (.A1(_054_),
    .A2(_059_),
    .ZN(_060_));
 BUF_X4 _349_ (.A(_060_),
    .Z(_061_));
 CLKBUF_X2 _350_ (.A(\state[2] ),
    .Z(_062_));
 CLKBUF_X3 _351_ (.A(_062_),
    .Z(_063_));
 BUF_X2 _352_ (.A(\iter[3] ),
    .Z(_064_));
 BUF_X2 _353_ (.A(\iter[2] ),
    .Z(_065_));
 NOR2_X4 _354_ (.A1(_064_),
    .A2(_065_),
    .ZN(_066_));
 NAND2_X1 _355_ (.A1(_291_),
    .A2(_066_),
    .ZN(_067_));
 NAND2_X1 _356_ (.A1(_063_),
    .A2(_067_),
    .ZN(_068_));
 AOI21_X1 _357_ (.A(_053_),
    .B1(_061_),
    .B2(_068_),
    .ZN(_002_));
 AOI21_X1 _358_ (.A(_052_),
    .B1(\state[1] ),
    .B2(_055_),
    .ZN(_069_));
 INV_X2 _359_ (.A(_054_),
    .ZN(_070_));
 OAI21_X1 _360_ (.A(_069_),
    .B1(_059_),
    .B2(_070_),
    .ZN(_000_));
 NAND2_X1 _361_ (.A1(_056_),
    .A2(\state[1] ),
    .ZN(_071_));
 NAND3_X4 _362_ (.A1(_062_),
    .A2(_291_),
    .A3(_066_),
    .ZN(_072_));
 AOI21_X1 _363_ (.A(_053_),
    .B1(_071_),
    .B2(_072_),
    .ZN(_001_));
 INV_X1 _364_ (.A(_065_),
    .ZN(_073_));
 BUF_X2 _365_ (.A(\iter[0] ),
    .Z(_074_));
 BUF_X2 _366_ (.A(_292_),
    .Z(_075_));
 INV_X1 _367_ (.A(_075_),
    .ZN(_076_));
 BUF_X2 _368_ (.A(_293_),
    .Z(_077_));
 MUX2_X1 _369_ (.A(net6),
    .B(net2),
    .S(_077_),
    .Z(_078_));
 NOR3_X1 _370_ (.A1(_074_),
    .A2(_076_),
    .A3(_078_),
    .ZN(_079_));
 MUX2_X1 _371_ (.A(net8),
    .B(net4),
    .S(_077_),
    .Z(_080_));
 MUX2_X1 _372_ (.A(net7),
    .B(net3),
    .S(_077_),
    .Z(_081_));
 MUX2_X1 _373_ (.A(_080_),
    .B(_081_),
    .S(_074_),
    .Z(_082_));
 MUX2_X1 _374_ (.A(net5),
    .B(net1),
    .S(_077_),
    .Z(_083_));
 NAND2_X1 _375_ (.A1(_074_),
    .A2(_075_),
    .ZN(_084_));
 OAI22_X1 _376_ (.A1(_075_),
    .A2(_082_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_085_));
 NOR4_X1 _377_ (.A1(_064_),
    .A2(_073_),
    .A3(_079_),
    .A4(_085_),
    .ZN(_086_));
 MUX2_X1 _378_ (.A(net8),
    .B(net6),
    .S(_075_),
    .Z(_087_));
 MUX2_X1 _379_ (.A(net7),
    .B(net5),
    .S(_075_),
    .Z(_088_));
 MUX2_X1 _380_ (.A(_087_),
    .B(_088_),
    .S(_074_),
    .Z(_089_));
 NAND3_X1 _381_ (.A1(_064_),
    .A2(_077_),
    .A3(_089_),
    .ZN(_090_));
 MUX2_X1 _382_ (.A(net4),
    .B(net2),
    .S(_075_),
    .Z(_091_));
 MUX2_X1 _383_ (.A(net3),
    .B(net1),
    .S(_075_),
    .Z(_092_));
 MUX2_X1 _384_ (.A(_091_),
    .B(_092_),
    .S(_074_),
    .Z(_093_));
 INV_X1 _385_ (.A(_093_),
    .ZN(_094_));
 OAI21_X1 _386_ (.A(_090_),
    .B1(_094_),
    .B2(_077_),
    .ZN(_095_));
 NOR3_X1 _387_ (.A1(_065_),
    .A2(_074_),
    .A3(\iter[1] ),
    .ZN(_096_));
 XOR2_X2 _388_ (.A(_064_),
    .B(_096_),
    .Z(_097_));
 NOR2_X1 _389_ (.A1(_065_),
    .A2(_097_),
    .ZN(_098_));
 AOI21_X2 _390_ (.A(_086_),
    .B1(_095_),
    .B2(_098_),
    .ZN(_299_));
 INV_X1 _391_ (.A(_299_),
    .ZN(_296_));
 BUF_X2 _392_ (.A(_051_),
    .Z(_099_));
 BUF_X2 _393_ (.A(_099_),
    .Z(_100_));
 INV_X2 _394_ (.A(_003_),
    .ZN(_101_));
 NAND2_X1 _395_ (.A1(_057_),
    .A2(_058_),
    .ZN(_102_));
 NAND2_X2 _396_ (.A1(_055_),
    .A2(_102_),
    .ZN(_103_));
 NOR2_X1 _397_ (.A1(_101_),
    .A2(_103_),
    .ZN(_104_));
 OAI21_X1 _398_ (.A(_072_),
    .B1(_063_),
    .B2(_070_),
    .ZN(_105_));
 MUX2_X1 _399_ (.A(net17),
    .B(_104_),
    .S(_105_),
    .Z(_106_));
 AND2_X1 _400_ (.A1(_100_),
    .A2(_106_),
    .ZN(_004_));
 MUX2_X1 _401_ (.A(net9),
    .B(\div_reg[0] ),
    .S(_061_),
    .Z(_107_));
 AND2_X1 _402_ (.A1(_100_),
    .A2(_107_),
    .ZN(_005_));
 MUX2_X1 _403_ (.A(net10),
    .B(\div_reg[1] ),
    .S(_061_),
    .Z(_108_));
 AND2_X1 _404_ (.A1(_100_),
    .A2(_108_),
    .ZN(_006_));
 NAND2_X1 _405_ (.A1(\div_reg[2] ),
    .A2(_061_),
    .ZN(_109_));
 NAND3_X1 _406_ (.A1(_055_),
    .A2(net11),
    .A3(_054_),
    .ZN(_110_));
 AOI21_X1 _407_ (.A(_053_),
    .B1(_109_),
    .B2(_110_),
    .ZN(_007_));
 MUX2_X1 _408_ (.A(net12),
    .B(\div_reg[3] ),
    .S(_061_),
    .Z(_111_));
 AND2_X1 _409_ (.A1(_100_),
    .A2(_111_),
    .ZN(_008_));
 MUX2_X1 _410_ (.A(net13),
    .B(\div_reg[4] ),
    .S(_061_),
    .Z(_112_));
 AND2_X1 _411_ (.A1(_100_),
    .A2(_112_),
    .ZN(_009_));
 MUX2_X1 _412_ (.A(net14),
    .B(\div_reg[5] ),
    .S(_061_),
    .Z(_113_));
 AND2_X1 _413_ (.A1(_100_),
    .A2(_113_),
    .ZN(_010_));
 MUX2_X1 _414_ (.A(net15),
    .B(\div_reg[6] ),
    .S(_061_),
    .Z(_114_));
 AND2_X1 _415_ (.A1(_100_),
    .A2(_114_),
    .ZN(_011_));
 MUX2_X1 _416_ (.A(net16),
    .B(\div_reg[7] ),
    .S(_061_),
    .Z(_115_));
 AND2_X1 _417_ (.A1(_100_),
    .A2(_115_),
    .ZN(_012_));
 NAND2_X1 _418_ (.A1(_070_),
    .A2(net18),
    .ZN(_116_));
 NAND4_X1 _419_ (.A1(_055_),
    .A2(_054_),
    .A3(_057_),
    .A4(_058_),
    .ZN(_117_));
 AOI21_X1 _420_ (.A(_053_),
    .B1(_116_),
    .B2(_117_),
    .ZN(_013_));
 AOI21_X2 _421_ (.A(_068_),
    .B1(_103_),
    .B2(_054_),
    .ZN(_118_));
 OR2_X2 _422_ (.A1(_054_),
    .A2(_062_),
    .ZN(_119_));
 OAI211_X4 _423_ (.A(_072_),
    .B(_119_),
    .C1(_070_),
    .C2(_059_),
    .ZN(_120_));
 MUX2_X1 _424_ (.A(_118_),
    .B(_120_),
    .S(_074_),
    .Z(_121_));
 AND2_X1 _425_ (.A1(_100_),
    .A2(_121_),
    .ZN(_014_));
 BUF_X4 _426_ (.A(_120_),
    .Z(_122_));
 AOI22_X1 _427_ (.A1(\iter[1] ),
    .A2(_122_),
    .B1(_118_),
    .B2(_076_),
    .ZN(_123_));
 NOR2_X1 _428_ (.A1(_053_),
    .A2(_123_),
    .ZN(_015_));
 XOR2_X1 _429_ (.A(_065_),
    .B(_077_),
    .Z(_124_));
 AOI22_X1 _430_ (.A1(_065_),
    .A2(_122_),
    .B1(_118_),
    .B2(_124_),
    .ZN(_125_));
 NOR2_X1 _431_ (.A1(_053_),
    .A2(_125_),
    .ZN(_016_));
 NAND2_X1 _432_ (.A1(_072_),
    .A2(_119_),
    .ZN(_126_));
 AOI21_X4 _433_ (.A(_126_),
    .B1(_103_),
    .B2(_054_),
    .ZN(_127_));
 NOR2_X1 _434_ (.A1(_064_),
    .A2(_127_),
    .ZN(_128_));
 NOR3_X1 _435_ (.A1(_003_),
    .A2(_097_),
    .A3(_120_),
    .ZN(_129_));
 NOR3_X1 _436_ (.A1(_053_),
    .A2(_128_),
    .A3(_129_),
    .ZN(_017_));
 INV_X2 _437_ (.A(_320_),
    .ZN(_130_));
 BUF_X2 _438_ (.A(_323_),
    .Z(_131_));
 INV_X2 _439_ (.A(_131_),
    .ZN(_132_));
 BUF_X4 _440_ (.A(_329_),
    .Z(_133_));
 INV_X4 _441_ (.A(_133_),
    .ZN(_134_));
 INV_X1 _442_ (.A(_335_),
    .ZN(_135_));
 NOR4_X2 _443_ (.A1(_130_),
    .A2(_132_),
    .A3(_134_),
    .A4(_135_),
    .ZN(_136_));
 BUF_X4 _444_ (.A(_308_),
    .Z(_137_));
 BUF_X4 _445_ (.A(_314_),
    .Z(_138_));
 AND2_X1 _446_ (.A1(_137_),
    .A2(_138_),
    .ZN(_139_));
 AND4_X1 _447_ (.A1(_303_),
    .A2(_298_),
    .A3(_136_),
    .A4(_139_),
    .ZN(_140_));
 INV_X1 _448_ (.A(_310_),
    .ZN(_141_));
 NAND3_X1 _449_ (.A1(_303_),
    .A2(_137_),
    .A3(_138_),
    .ZN(_142_));
 AOI21_X1 _450_ (.A(_316_),
    .B1(_138_),
    .B2(_304_),
    .ZN(_143_));
 INV_X1 _451_ (.A(_137_),
    .ZN(_144_));
 OAI221_X2 _452_ (.A(_141_),
    .B1(_142_),
    .B2(_297_),
    .C1(_143_),
    .C2(_144_),
    .ZN(_145_));
 INV_X1 _453_ (.A(_325_),
    .ZN(_146_));
 AOI21_X1 _454_ (.A(_331_),
    .B1(_133_),
    .B2(_337_),
    .ZN(_147_));
 OAI21_X1 _455_ (.A(_146_),
    .B1(_132_),
    .B2(_147_),
    .ZN(_148_));
 AOI221_X2 _456_ (.A(_319_),
    .B1(_136_),
    .B2(_145_),
    .C1(_148_),
    .C2(_320_),
    .ZN(_149_));
 OR2_X1 _457_ (.A1(_140_),
    .A2(_149_),
    .ZN(_150_));
 BUF_X8 _458_ (.A(_150_),
    .Z(_151_));
 AOI22_X1 _459_ (.A1(\quot[0] ),
    .A2(_122_),
    .B1(_118_),
    .B2(_151_),
    .ZN(_152_));
 NOR2_X1 _460_ (.A1(_053_),
    .A2(_152_),
    .ZN(_018_));
 NAND2_X1 _461_ (.A1(\quot[1] ),
    .A2(_122_),
    .ZN(_153_));
 NAND3_X1 _462_ (.A1(_063_),
    .A2(\quot[0] ),
    .A3(_127_),
    .ZN(_154_));
 AOI21_X1 _463_ (.A(_053_),
    .B1(_153_),
    .B2(_154_),
    .ZN(_019_));
 NAND2_X1 _464_ (.A1(\quot[2] ),
    .A2(_122_),
    .ZN(_155_));
 NAND3_X1 _465_ (.A1(_063_),
    .A2(\quot[1] ),
    .A3(_127_),
    .ZN(_156_));
 AOI21_X1 _466_ (.A(_053_),
    .B1(_155_),
    .B2(_156_),
    .ZN(_020_));
 NAND2_X1 _467_ (.A1(\quot[3] ),
    .A2(_122_),
    .ZN(_157_));
 NAND3_X1 _468_ (.A1(_063_),
    .A2(\quot[2] ),
    .A3(_127_),
    .ZN(_158_));
 AOI21_X1 _469_ (.A(_052_),
    .B1(_157_),
    .B2(_158_),
    .ZN(_021_));
 NAND2_X1 _470_ (.A1(\quot[4] ),
    .A2(_122_),
    .ZN(_159_));
 NAND3_X1 _471_ (.A1(_063_),
    .A2(\quot[3] ),
    .A3(_127_),
    .ZN(_160_));
 AOI21_X1 _472_ (.A(_052_),
    .B1(_159_),
    .B2(_160_),
    .ZN(_022_));
 NAND2_X1 _473_ (.A1(\quot[5] ),
    .A2(_122_),
    .ZN(_161_));
 NAND3_X1 _474_ (.A1(_063_),
    .A2(\quot[4] ),
    .A3(_127_),
    .ZN(_162_));
 AOI21_X1 _475_ (.A(_052_),
    .B1(_161_),
    .B2(_162_),
    .ZN(_023_));
 NAND2_X1 _476_ (.A1(\quot[6] ),
    .A2(_122_),
    .ZN(_163_));
 NAND3_X1 _477_ (.A1(_063_),
    .A2(\quot[5] ),
    .A3(_127_),
    .ZN(_164_));
 AOI21_X1 _478_ (.A(_052_),
    .B1(_163_),
    .B2(_164_),
    .ZN(_024_));
 NAND2_X1 _479_ (.A1(\quot[7] ),
    .A2(_122_),
    .ZN(_165_));
 NAND3_X1 _480_ (.A1(_063_),
    .A2(\quot[6] ),
    .A3(_127_),
    .ZN(_166_));
 AOI21_X1 _481_ (.A(_052_),
    .B1(_165_),
    .B2(_166_),
    .ZN(_025_));
 NAND3_X4 _482_ (.A1(_101_),
    .A2(_291_),
    .A3(_066_),
    .ZN(_167_));
 CLKBUF_X3 _483_ (.A(_167_),
    .Z(_168_));
 MUX2_X1 _484_ (.A(\quot[0] ),
    .B(net19),
    .S(_168_),
    .Z(_169_));
 AND2_X1 _485_ (.A1(_100_),
    .A2(_169_),
    .ZN(_026_));
 BUF_X2 _486_ (.A(_099_),
    .Z(_170_));
 MUX2_X1 _487_ (.A(\quot[1] ),
    .B(net20),
    .S(_168_),
    .Z(_171_));
 AND2_X1 _488_ (.A1(_170_),
    .A2(_171_),
    .ZN(_027_));
 MUX2_X1 _489_ (.A(\quot[2] ),
    .B(net21),
    .S(_168_),
    .Z(_172_));
 AND2_X1 _490_ (.A1(_170_),
    .A2(_172_),
    .ZN(_028_));
 MUX2_X1 _491_ (.A(\quot[3] ),
    .B(net22),
    .S(_168_),
    .Z(_173_));
 AND2_X1 _492_ (.A1(_170_),
    .A2(_173_),
    .ZN(_029_));
 MUX2_X1 _493_ (.A(\quot[4] ),
    .B(net23),
    .S(_168_),
    .Z(_174_));
 AND2_X1 _494_ (.A1(_170_),
    .A2(_174_),
    .ZN(_030_));
 MUX2_X1 _495_ (.A(\quot[5] ),
    .B(net24),
    .S(_168_),
    .Z(_175_));
 AND2_X1 _496_ (.A1(_170_),
    .A2(_175_),
    .ZN(_031_));
 MUX2_X1 _497_ (.A(\quot[6] ),
    .B(net25),
    .S(_168_),
    .Z(_176_));
 AND2_X1 _498_ (.A1(_170_),
    .A2(_176_),
    .ZN(_032_));
 MUX2_X1 _499_ (.A(\quot[7] ),
    .B(net26),
    .S(_168_),
    .Z(_177_));
 AND2_X1 _500_ (.A1(_170_),
    .A2(_177_),
    .ZN(_033_));
 INV_X1 _501_ (.A(_298_),
    .ZN(_178_));
 NAND3_X2 _502_ (.A1(_051_),
    .A2(_101_),
    .A3(_072_),
    .ZN(_179_));
 NAND2_X1 _503_ (.A1(_070_),
    .A2(_062_),
    .ZN(_180_));
 AOI21_X4 _504_ (.A(_179_),
    .B1(_180_),
    .B2(_061_),
    .ZN(_181_));
 NAND3_X1 _505_ (.A1(_178_),
    .A2(_149_),
    .A3(_181_),
    .ZN(_182_));
 NOR2_X1 _506_ (.A1(_140_),
    .A2(_149_),
    .ZN(_183_));
 NAND2_X1 _507_ (.A1(_183_),
    .A2(_181_),
    .ZN(_184_));
 INV_X1 _508_ (.A(\rem[0] ),
    .ZN(_185_));
 NAND2_X2 _509_ (.A1(_099_),
    .A2(_120_),
    .ZN(_186_));
 OAI221_X1 _510_ (.A(_182_),
    .B1(_184_),
    .B2(_299_),
    .C1(_185_),
    .C2(_186_),
    .ZN(_034_));
 NAND3_X1 _511_ (.A1(_288_),
    .A2(_151_),
    .A3(_181_),
    .ZN(_187_));
 NAND2_X1 _512_ (.A1(\rem[0] ),
    .A2(_181_),
    .ZN(_188_));
 INV_X1 _513_ (.A(\rem[1] ),
    .ZN(_189_));
 OAI221_X1 _514_ (.A(_187_),
    .B1(_188_),
    .B2(_151_),
    .C1(_186_),
    .C2(_189_),
    .ZN(_035_));
 INV_X1 _515_ (.A(\rem[2] ),
    .ZN(_190_));
 AND2_X1 _516_ (.A1(_060_),
    .A2(_180_),
    .ZN(_191_));
 OR2_X2 _517_ (.A1(_191_),
    .A2(_179_),
    .ZN(_192_));
 XOR2_X1 _518_ (.A(_287_),
    .B(_138_),
    .Z(_193_));
 MUX2_X1 _519_ (.A(_189_),
    .B(_193_),
    .S(_151_),
    .Z(_194_));
 OAI22_X1 _520_ (.A1(_190_),
    .A2(_186_),
    .B1(_192_),
    .B2(_194_),
    .ZN(_036_));
 INV_X1 _521_ (.A(\rem[3] ),
    .ZN(_195_));
 INV_X1 _522_ (.A(_313_),
    .ZN(_196_));
 INV_X1 _523_ (.A(_286_),
    .ZN(_197_));
 AOI21_X2 _524_ (.A(_302_),
    .B1(_197_),
    .B2(_303_),
    .ZN(_198_));
 INV_X1 _525_ (.A(_138_),
    .ZN(_199_));
 OAI21_X1 _526_ (.A(_196_),
    .B1(_198_),
    .B2(_199_),
    .ZN(_200_));
 XNOR2_X1 _527_ (.A(_137_),
    .B(_200_),
    .ZN(_201_));
 MUX2_X1 _528_ (.A(_190_),
    .B(_201_),
    .S(_151_),
    .Z(_202_));
 OAI22_X1 _529_ (.A1(_195_),
    .A2(_186_),
    .B1(_192_),
    .B2(_202_),
    .ZN(_037_));
 INV_X1 _530_ (.A(\rem[4] ),
    .ZN(_203_));
 OR2_X1 _531_ (.A1(_307_),
    .A2(_313_),
    .ZN(_204_));
 INV_X1 _532_ (.A(_287_),
    .ZN(_205_));
 AOI21_X1 _533_ (.A(_204_),
    .B1(_138_),
    .B2(_205_),
    .ZN(_206_));
 NOR2_X1 _534_ (.A1(_137_),
    .A2(_307_),
    .ZN(_207_));
 NOR2_X1 _535_ (.A1(_206_),
    .A2(_207_),
    .ZN(_208_));
 XNOR2_X1 _536_ (.A(_335_),
    .B(_208_),
    .ZN(_209_));
 MUX2_X1 _537_ (.A(_195_),
    .B(_209_),
    .S(_151_),
    .Z(_210_));
 OAI22_X1 _538_ (.A1(_203_),
    .A2(_186_),
    .B1(_192_),
    .B2(_210_),
    .ZN(_038_));
 AND2_X1 _539_ (.A1(_099_),
    .A2(_120_),
    .ZN(_211_));
 NAND2_X1 _540_ (.A1(\rem[5] ),
    .A2(_211_),
    .ZN(_212_));
 INV_X1 _541_ (.A(_334_),
    .ZN(_213_));
 NAND2_X1 _542_ (.A1(_335_),
    .A2(_139_),
    .ZN(_214_));
 AOI21_X1 _543_ (.A(_307_),
    .B1(_313_),
    .B2(_137_),
    .ZN(_215_));
 OAI221_X2 _544_ (.A(_213_),
    .B1(_198_),
    .B2(_214_),
    .C1(_215_),
    .C2(_135_),
    .ZN(_216_));
 XNOR2_X1 _545_ (.A(_133_),
    .B(_216_),
    .ZN(_217_));
 MUX2_X1 _546_ (.A(_203_),
    .B(_217_),
    .S(_151_),
    .Z(_218_));
 OAI21_X1 _547_ (.A(_212_),
    .B1(_218_),
    .B2(_192_),
    .ZN(_039_));
 NAND3_X1 _548_ (.A1(\rem[5] ),
    .A2(_183_),
    .A3(_181_),
    .ZN(_219_));
 CLKBUF_X2 _549_ (.A(_328_),
    .Z(_220_));
 NOR3_X1 _550_ (.A1(_132_),
    .A2(_220_),
    .A3(_334_),
    .ZN(_221_));
 NOR2_X1 _551_ (.A1(_131_),
    .A2(_134_),
    .ZN(_222_));
 NOR3_X1 _552_ (.A1(_135_),
    .A2(_206_),
    .A3(_207_),
    .ZN(_223_));
 MUX2_X1 _553_ (.A(_221_),
    .B(_222_),
    .S(_223_),
    .Z(_224_));
 NOR3_X1 _554_ (.A1(_132_),
    .A2(_133_),
    .A3(_220_),
    .ZN(_225_));
 AOI21_X1 _555_ (.A(_225_),
    .B1(_222_),
    .B2(_334_),
    .ZN(_226_));
 INV_X1 _556_ (.A(_220_),
    .ZN(_227_));
 OAI21_X1 _557_ (.A(_226_),
    .B1(_227_),
    .B2(_131_),
    .ZN(_228_));
 OAI21_X1 _558_ (.A(_151_),
    .B1(_224_),
    .B2(_228_),
    .ZN(_229_));
 INV_X1 _559_ (.A(\rem[6] ),
    .ZN(_230_));
 OAI221_X1 _560_ (.A(_219_),
    .B1(_229_),
    .B2(_192_),
    .C1(_230_),
    .C2(_186_),
    .ZN(_040_));
 INV_X1 _561_ (.A(\rem[7] ),
    .ZN(_231_));
 NOR2_X1 _562_ (.A1(\rem[6] ),
    .A2(_151_),
    .ZN(_232_));
 AND4_X1 _563_ (.A1(_130_),
    .A2(_131_),
    .A3(_133_),
    .A4(_216_),
    .ZN(_233_));
 NOR4_X1 _564_ (.A1(_130_),
    .A2(_322_),
    .A3(_220_),
    .A4(_216_),
    .ZN(_234_));
 OR4_X1 _565_ (.A1(_130_),
    .A2(_133_),
    .A3(_322_),
    .A4(_220_),
    .ZN(_235_));
 NAND3_X1 _566_ (.A1(_130_),
    .A2(_131_),
    .A3(_220_),
    .ZN(_236_));
 NOR3_X1 _567_ (.A1(_130_),
    .A2(_131_),
    .A3(_322_),
    .ZN(_237_));
 AOI21_X1 _568_ (.A(_237_),
    .B1(_322_),
    .B2(_130_),
    .ZN(_238_));
 NAND3_X1 _569_ (.A1(_235_),
    .A2(_236_),
    .A3(_238_),
    .ZN(_239_));
 NOR4_X1 _570_ (.A1(_183_),
    .A2(_233_),
    .A3(_234_),
    .A4(_239_),
    .ZN(_240_));
 OAI33_X1 _571_ (.A1(_052_),
    .A2(_231_),
    .A3(_127_),
    .B1(_192_),
    .B2(_232_),
    .B3(_240_),
    .ZN(_041_));
 MUX2_X1 _572_ (.A(\rem[0] ),
    .B(net27),
    .S(_168_),
    .Z(_241_));
 AND2_X1 _573_ (.A1(_170_),
    .A2(_241_),
    .ZN(_042_));
 MUX2_X1 _574_ (.A(\rem[1] ),
    .B(net28),
    .S(_168_),
    .Z(_242_));
 AND2_X1 _575_ (.A1(_170_),
    .A2(_242_),
    .ZN(_043_));
 MUX2_X1 _576_ (.A(\rem[2] ),
    .B(net29),
    .S(_167_),
    .Z(_243_));
 AND2_X1 _577_ (.A1(_170_),
    .A2(_243_),
    .ZN(_044_));
 MUX2_X1 _578_ (.A(\rem[3] ),
    .B(net30),
    .S(_167_),
    .Z(_244_));
 AND2_X1 _579_ (.A1(_099_),
    .A2(_244_),
    .ZN(_045_));
 MUX2_X1 _580_ (.A(\rem[4] ),
    .B(net31),
    .S(_167_),
    .Z(_245_));
 AND2_X1 _581_ (.A1(_099_),
    .A2(_245_),
    .ZN(_046_));
 MUX2_X1 _582_ (.A(\rem[5] ),
    .B(net32),
    .S(_167_),
    .Z(_246_));
 AND2_X1 _583_ (.A1(_099_),
    .A2(_246_),
    .ZN(_047_));
 MUX2_X1 _584_ (.A(\rem[6] ),
    .B(net33),
    .S(_167_),
    .Z(_247_));
 AND2_X1 _585_ (.A1(_099_),
    .A2(_247_),
    .ZN(_048_));
 MUX2_X1 _586_ (.A(\rem[7] ),
    .B(net34),
    .S(_167_),
    .Z(_248_));
 AND2_X1 _587_ (.A1(_099_),
    .A2(_248_),
    .ZN(_049_));
 OAI21_X1 _588_ (.A(_071_),
    .B1(_119_),
    .B2(\state[1] ),
    .ZN(_249_));
 NOR2_X1 _589_ (.A1(_067_),
    .A2(_249_),
    .ZN(_250_));
 OAI221_X1 _590_ (.A(_099_),
    .B1(_063_),
    .B2(_249_),
    .C1(_250_),
    .C2(net35),
    .ZN(_251_));
 INV_X1 _591_ (.A(_251_),
    .ZN(_050_));
 FA_X1 _592_ (.A(\div_reg[1] ),
    .B(_285_),
    .CI(_286_),
    .CO(_287_),
    .S(_288_));
 HA_X1 _593_ (.A(_289_),
    .B(_290_),
    .CO(_291_),
    .S(_292_));
 HA_X1 _594_ (.A(_289_),
    .B(_290_),
    .CO(_293_),
    .S(_294_));
 HA_X1 _595_ (.A(_295_),
    .B(_296_),
    .CO(_297_),
    .S(_298_));
 HA_X1 _596_ (.A(\div_reg[0] ),
    .B(_299_),
    .CO(_286_),
    .S(_300_));
 HA_X1 _597_ (.A(_301_),
    .B(\rem[0] ),
    .CO(_302_),
    .S(_303_));
 HA_X1 _598_ (.A(\div_reg[1] ),
    .B(_285_),
    .CO(_304_),
    .S(_305_));
 HA_X1 _599_ (.A(_306_),
    .B(\rem[2] ),
    .CO(_307_),
    .S(_308_));
 HA_X1 _600_ (.A(\div_reg[3] ),
    .B(_309_),
    .CO(_310_),
    .S(_311_));
 HA_X1 _601_ (.A(_312_),
    .B(\rem[1] ),
    .CO(_313_),
    .S(_314_));
 HA_X1 _602_ (.A(\div_reg[2] ),
    .B(_315_),
    .CO(_316_),
    .S(_317_));
 HA_X1 _603_ (.A(\div_reg[7] ),
    .B(_318_),
    .CO(_319_),
    .S(_320_));
 HA_X1 _604_ (.A(_321_),
    .B(\rem[5] ),
    .CO(_322_),
    .S(_323_));
 HA_X1 _605_ (.A(\div_reg[6] ),
    .B(_324_),
    .CO(_325_),
    .S(_326_));
 HA_X1 _606_ (.A(_327_),
    .B(\rem[4] ),
    .CO(_328_),
    .S(_329_));
 HA_X1 _607_ (.A(\div_reg[5] ),
    .B(_330_),
    .CO(_331_),
    .S(_332_));
 HA_X1 _608_ (.A(_333_),
    .B(\rem[3] ),
    .CO(_334_),
    .S(_335_));
 HA_X1 _609_ (.A(\div_reg[4] ),
    .B(_336_),
    .CO(_337_),
    .S(_338_));
 DFF_X1 \busy$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_281_));
 DFF_X1 \div_reg[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\div_reg[0] ),
    .QN(_295_));
 DFF_X2 \div_reg[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\div_reg[1] ),
    .QN(_301_));
 DFF_X1 \div_reg[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\div_reg[2] ),
    .QN(_312_));
 DFF_X1 \div_reg[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\div_reg[3] ),
    .QN(_306_));
 DFF_X1 \div_reg[4]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\div_reg[4] ),
    .QN(_333_));
 DFF_X1 \div_reg[5]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\div_reg[5] ),
    .QN(_327_));
 DFF_X1 \div_reg[6]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\div_reg[6] ),
    .QN(_321_));
 DFF_X1 \div_reg[7]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\div_reg[7] ),
    .QN(_280_));
 DFF_X1 \error$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net18),
    .QN(_279_));
 DFF_X1 \iter[0]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\iter[0] ),
    .QN(_289_));
 DFF_X1 \iter[1]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\iter[1] ),
    .QN(_290_));
 DFF_X1 \iter[2]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\iter[2] ),
    .QN(_278_));
 DFF_X1 \iter[3]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\iter[3] ),
    .QN(_277_));
 DFF_X1 \quot[0]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\quot[0] ),
    .QN(_276_));
 DFF_X1 \quot[1]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\quot[1] ),
    .QN(_275_));
 DFF_X1 \quot[2]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\quot[2] ),
    .QN(_274_));
 DFF_X1 \quot[3]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\quot[3] ),
    .QN(_273_));
 DFF_X1 \quot[4]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\quot[4] ),
    .QN(_272_));
 DFF_X1 \quot[5]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\quot[5] ),
    .QN(_271_));
 DFF_X1 \quot[6]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\quot[6] ),
    .QN(_270_));
 DFF_X1 \quot[7]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\quot[7] ),
    .QN(_269_));
 DFF_X1 \quotient[0]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net19),
    .QN(_268_));
 DFF_X1 \quotient[1]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net20),
    .QN(_267_));
 DFF_X1 \quotient[2]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net21),
    .QN(_266_));
 DFF_X1 \quotient[3]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net22),
    .QN(_265_));
 DFF_X1 \quotient[4]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net23),
    .QN(_264_));
 DFF_X1 \quotient[5]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net24),
    .QN(_263_));
 DFF_X1 \quotient[6]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net25),
    .QN(_262_));
 DFF_X1 \quotient[7]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net26),
    .QN(_261_));
 DFF_X2 \rem[0]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\rem[0] ),
    .QN(_285_));
 DFF_X1 \rem[1]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\rem[1] ),
    .QN(_315_));
 DFF_X1 \rem[2]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rem[2] ),
    .QN(_309_));
 DFF_X1 \rem[3]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rem[3] ),
    .QN(_336_));
 DFF_X1 \rem[4]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rem[4] ),
    .QN(_330_));
 DFF_X2 \rem[5]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rem[5] ),
    .QN(_324_));
 DFF_X1 \rem[6]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rem[6] ),
    .QN(_318_));
 DFF_X1 \rem[7]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rem[7] ),
    .QN(_260_));
 DFF_X1 \remainder[0]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net27),
    .QN(_259_));
 DFF_X1 \remainder[1]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net28),
    .QN(_258_));
 DFF_X1 \remainder[2]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net29),
    .QN(_257_));
 DFF_X1 \remainder[3]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net30),
    .QN(_256_));
 DFF_X1 \remainder[4]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net31),
    .QN(_255_));
 DFF_X1 \remainder[5]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net32),
    .QN(_254_));
 DFF_X1 \remainder[6]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net33),
    .QN(_253_));
 DFF_X1 \remainder[7]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net34),
    .QN(_282_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[0] ),
    .QN(_283_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\state[1] ),
    .QN(_284_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[2] ),
    .QN(_003_));
 DFF_X1 \valid$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net35),
    .QN(_252_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 BUF_X1 input1 (.A(dividend[0]),
    .Z(net1));
 BUF_X1 input2 (.A(dividend[1]),
    .Z(net2));
 BUF_X1 input3 (.A(dividend[2]),
    .Z(net3));
 BUF_X1 input4 (.A(dividend[3]),
    .Z(net4));
 BUF_X1 input5 (.A(dividend[4]),
    .Z(net5));
 BUF_X1 input6 (.A(dividend[5]),
    .Z(net6));
 BUF_X1 input7 (.A(dividend[6]),
    .Z(net7));
 BUF_X1 input8 (.A(dividend[7]),
    .Z(net8));
 BUF_X1 input9 (.A(divisor[0]),
    .Z(net9));
 BUF_X1 input10 (.A(divisor[1]),
    .Z(net10));
 BUF_X1 input11 (.A(divisor[2]),
    .Z(net11));
 BUF_X1 input12 (.A(divisor[3]),
    .Z(net12));
 BUF_X1 input13 (.A(divisor[4]),
    .Z(net13));
 BUF_X1 input14 (.A(divisor[5]),
    .Z(net14));
 BUF_X1 input15 (.A(divisor[6]),
    .Z(net15));
 BUF_X1 input16 (.A(divisor[7]),
    .Z(net16));
 BUF_X1 output17 (.A(net17),
    .Z(busy));
 BUF_X1 output18 (.A(net18),
    .Z(error));
 BUF_X1 output19 (.A(net19),
    .Z(quotient[0]));
 BUF_X1 output20 (.A(net20),
    .Z(quotient[1]));
 BUF_X1 output21 (.A(net21),
    .Z(quotient[2]));
 BUF_X1 output22 (.A(net22),
    .Z(quotient[3]));
 BUF_X1 output23 (.A(net23),
    .Z(quotient[4]));
 BUF_X1 output24 (.A(net24),
    .Z(quotient[5]));
 BUF_X1 output25 (.A(net25),
    .Z(quotient[6]));
 BUF_X1 output26 (.A(net26),
    .Z(quotient[7]));
 BUF_X1 output27 (.A(net27),
    .Z(remainder[0]));
 BUF_X1 output28 (.A(net28),
    .Z(remainder[1]));
 BUF_X1 output29 (.A(net29),
    .Z(remainder[2]));
 BUF_X1 output30 (.A(net30),
    .Z(remainder[3]));
 BUF_X1 output31 (.A(net31),
    .Z(remainder[4]));
 BUF_X1 output32 (.A(net32),
    .Z(remainder[5]));
 BUF_X1 output33 (.A(net33),
    .Z(remainder[6]));
 BUF_X1 output34 (.A(net34),
    .Z(remainder[7]));
 BUF_X1 output35 (.A(net35),
    .Z(valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X4 clkload1 (.A(clknet_2_1__leaf_clk));
 INV_X1 clkload2 (.A(clknet_2_2__leaf_clk));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X1 FILLER_0_17 ();
 FILLCELL_X2 FILLER_0_24 ();
 FILLCELL_X1 FILLER_0_26 ();
 FILLCELL_X16 FILLER_0_30 ();
 FILLCELL_X2 FILLER_0_46 ();
 FILLCELL_X1 FILLER_0_48 ();
 FILLCELL_X4 FILLER_0_55 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_89 ();
 FILLCELL_X32 FILLER_0_100 ();
 FILLCELL_X32 FILLER_0_132 ();
 FILLCELL_X8 FILLER_0_164 ();
 FILLCELL_X4 FILLER_0_172 ();
 FILLCELL_X1 FILLER_0_176 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X8 FILLER_1_27 ();
 FILLCELL_X1 FILLER_1_35 ();
 FILLCELL_X4 FILLER_1_54 ();
 FILLCELL_X2 FILLER_1_69 ();
 FILLCELL_X1 FILLER_1_71 ();
 FILLCELL_X2 FILLER_1_96 ();
 FILLCELL_X1 FILLER_1_98 ();
 FILLCELL_X2 FILLER_1_101 ();
 FILLCELL_X1 FILLER_1_103 ();
 FILLCELL_X32 FILLER_1_114 ();
 FILLCELL_X16 FILLER_1_146 ();
 FILLCELL_X8 FILLER_1_162 ();
 FILLCELL_X4 FILLER_1_170 ();
 FILLCELL_X2 FILLER_1_174 ();
 FILLCELL_X1 FILLER_1_176 ();
 FILLCELL_X2 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_3 ();
 FILLCELL_X4 FILLER_2_7 ();
 FILLCELL_X2 FILLER_2_11 ();
 FILLCELL_X8 FILLER_2_34 ();
 FILLCELL_X2 FILLER_2_42 ();
 FILLCELL_X1 FILLER_2_44 ();
 FILLCELL_X4 FILLER_2_75 ();
 FILLCELL_X8 FILLER_2_83 ();
 FILLCELL_X2 FILLER_2_91 ();
 FILLCELL_X32 FILLER_2_110 ();
 FILLCELL_X32 FILLER_2_142 ();
 FILLCELL_X2 FILLER_2_174 ();
 FILLCELL_X1 FILLER_2_176 ();
 FILLCELL_X4 FILLER_3_1 ();
 FILLCELL_X2 FILLER_3_12 ();
 FILLCELL_X1 FILLER_3_14 ();
 FILLCELL_X1 FILLER_3_22 ();
 FILLCELL_X4 FILLER_3_30 ();
 FILLCELL_X1 FILLER_3_34 ();
 FILLCELL_X4 FILLER_3_37 ();
 FILLCELL_X8 FILLER_3_58 ();
 FILLCELL_X1 FILLER_3_66 ();
 FILLCELL_X8 FILLER_3_87 ();
 FILLCELL_X1 FILLER_3_95 ();
 FILLCELL_X2 FILLER_3_102 ();
 FILLCELL_X32 FILLER_3_119 ();
 FILLCELL_X16 FILLER_3_151 ();
 FILLCELL_X8 FILLER_3_167 ();
 FILLCELL_X2 FILLER_3_175 ();
 FILLCELL_X1 FILLER_4_24 ();
 FILLCELL_X1 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_42 ();
 FILLCELL_X2 FILLER_4_46 ();
 FILLCELL_X1 FILLER_4_58 ();
 FILLCELL_X4 FILLER_4_75 ();
 FILLCELL_X2 FILLER_4_79 ();
 FILLCELL_X2 FILLER_4_83 ();
 FILLCELL_X1 FILLER_4_92 ();
 FILLCELL_X1 FILLER_4_97 ();
 FILLCELL_X1 FILLER_4_112 ();
 FILLCELL_X8 FILLER_4_150 ();
 FILLCELL_X8 FILLER_4_165 ();
 FILLCELL_X4 FILLER_4_173 ();
 FILLCELL_X2 FILLER_5_18 ();
 FILLCELL_X2 FILLER_5_26 ();
 FILLCELL_X1 FILLER_5_28 ();
 FILLCELL_X1 FILLER_5_36 ();
 FILLCELL_X8 FILLER_5_47 ();
 FILLCELL_X2 FILLER_5_55 ();
 FILLCELL_X1 FILLER_5_76 ();
 FILLCELL_X1 FILLER_5_81 ();
 FILLCELL_X1 FILLER_5_105 ();
 FILLCELL_X1 FILLER_5_108 ();
 FILLCELL_X1 FILLER_5_113 ();
 FILLCELL_X2 FILLER_5_118 ();
 FILLCELL_X1 FILLER_5_120 ();
 FILLCELL_X8 FILLER_5_136 ();
 FILLCELL_X1 FILLER_5_144 ();
 FILLCELL_X4 FILLER_5_155 ();
 FILLCELL_X2 FILLER_5_159 ();
 FILLCELL_X8 FILLER_5_165 ();
 FILLCELL_X4 FILLER_5_173 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_9 ();
 FILLCELL_X2 FILLER_6_13 ();
 FILLCELL_X1 FILLER_6_15 ();
 FILLCELL_X8 FILLER_6_22 ();
 FILLCELL_X2 FILLER_6_30 ();
 FILLCELL_X16 FILLER_6_46 ();
 FILLCELL_X8 FILLER_6_62 ();
 FILLCELL_X4 FILLER_6_70 ();
 FILLCELL_X1 FILLER_6_81 ();
 FILLCELL_X16 FILLER_6_90 ();
 FILLCELL_X4 FILLER_6_138 ();
 FILLCELL_X1 FILLER_6_142 ();
 FILLCELL_X16 FILLER_6_160 ();
 FILLCELL_X1 FILLER_6_176 ();
 FILLCELL_X1 FILLER_7_22 ();
 FILLCELL_X2 FILLER_7_27 ();
 FILLCELL_X1 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_44 ();
 FILLCELL_X4 FILLER_7_69 ();
 FILLCELL_X4 FILLER_7_83 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X1 FILLER_7_93 ();
 FILLCELL_X8 FILLER_7_100 ();
 FILLCELL_X2 FILLER_7_108 ();
 FILLCELL_X4 FILLER_7_124 ();
 FILLCELL_X2 FILLER_7_128 ();
 FILLCELL_X1 FILLER_7_130 ();
 FILLCELL_X8 FILLER_7_163 ();
 FILLCELL_X4 FILLER_7_171 ();
 FILLCELL_X2 FILLER_7_175 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_34 ();
 FILLCELL_X2 FILLER_8_42 ();
 FILLCELL_X2 FILLER_8_47 ();
 FILLCELL_X1 FILLER_8_49 ();
 FILLCELL_X8 FILLER_8_54 ();
 FILLCELL_X2 FILLER_8_62 ();
 FILLCELL_X1 FILLER_8_86 ();
 FILLCELL_X1 FILLER_8_91 ();
 FILLCELL_X1 FILLER_8_99 ();
 FILLCELL_X8 FILLER_8_123 ();
 FILLCELL_X4 FILLER_8_131 ();
 FILLCELL_X8 FILLER_8_167 ();
 FILLCELL_X2 FILLER_8_175 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_9 ();
 FILLCELL_X2 FILLER_9_13 ();
 FILLCELL_X1 FILLER_9_15 ();
 FILLCELL_X1 FILLER_9_53 ();
 FILLCELL_X2 FILLER_9_58 ();
 FILLCELL_X1 FILLER_9_60 ();
 FILLCELL_X1 FILLER_9_78 ();
 FILLCELL_X4 FILLER_9_88 ();
 FILLCELL_X2 FILLER_9_92 ();
 FILLCELL_X2 FILLER_9_105 ();
 FILLCELL_X2 FILLER_9_119 ();
 FILLCELL_X1 FILLER_9_121 ();
 FILLCELL_X2 FILLER_9_130 ();
 FILLCELL_X2 FILLER_9_134 ();
 FILLCELL_X1 FILLER_9_136 ();
 FILLCELL_X2 FILLER_9_141 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X1 FILLER_9_148 ();
 FILLCELL_X16 FILLER_9_151 ();
 FILLCELL_X8 FILLER_9_167 ();
 FILLCELL_X2 FILLER_9_175 ();
 FILLCELL_X4 FILLER_10_26 ();
 FILLCELL_X2 FILLER_10_30 ();
 FILLCELL_X4 FILLER_10_45 ();
 FILLCELL_X1 FILLER_10_49 ();
 FILLCELL_X32 FILLER_10_54 ();
 FILLCELL_X16 FILLER_10_86 ();
 FILLCELL_X4 FILLER_10_102 ();
 FILLCELL_X1 FILLER_10_106 ();
 FILLCELL_X2 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_141 ();
 FILLCELL_X4 FILLER_10_156 ();
 FILLCELL_X1 FILLER_10_160 ();
 FILLCELL_X4 FILLER_10_172 ();
 FILLCELL_X1 FILLER_10_176 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X4 FILLER_11_16 ();
 FILLCELL_X1 FILLER_11_20 ();
 FILLCELL_X1 FILLER_11_38 ();
 FILLCELL_X2 FILLER_11_43 ();
 FILLCELL_X2 FILLER_11_62 ();
 FILLCELL_X2 FILLER_11_71 ();
 FILLCELL_X1 FILLER_11_73 ();
 FILLCELL_X1 FILLER_11_78 ();
 FILLCELL_X8 FILLER_11_84 ();
 FILLCELL_X1 FILLER_11_109 ();
 FILLCELL_X2 FILLER_11_122 ();
 FILLCELL_X1 FILLER_11_124 ();
 FILLCELL_X16 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_145 ();
 FILLCELL_X1 FILLER_11_149 ();
 FILLCELL_X2 FILLER_11_157 ();
 FILLCELL_X1 FILLER_11_159 ();
 FILLCELL_X4 FILLER_12_18 ();
 FILLCELL_X4 FILLER_12_29 ();
 FILLCELL_X2 FILLER_12_36 ();
 FILLCELL_X2 FILLER_12_53 ();
 FILLCELL_X1 FILLER_12_55 ();
 FILLCELL_X4 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_70 ();
 FILLCELL_X2 FILLER_12_87 ();
 FILLCELL_X2 FILLER_12_94 ();
 FILLCELL_X1 FILLER_12_96 ();
 FILLCELL_X2 FILLER_12_107 ();
 FILLCELL_X4 FILLER_12_124 ();
 FILLCELL_X4 FILLER_12_142 ();
 FILLCELL_X2 FILLER_12_146 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_67 ();
 FILLCELL_X4 FILLER_13_81 ();
 FILLCELL_X2 FILLER_13_92 ();
 FILLCELL_X8 FILLER_13_101 ();
 FILLCELL_X2 FILLER_13_109 ();
 FILLCELL_X1 FILLER_13_122 ();
 FILLCELL_X4 FILLER_13_129 ();
 FILLCELL_X2 FILLER_13_133 ();
 FILLCELL_X4 FILLER_13_137 ();
 FILLCELL_X4 FILLER_13_158 ();
 FILLCELL_X2 FILLER_13_168 ();
 FILLCELL_X1 FILLER_13_170 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_17 ();
 FILLCELL_X2 FILLER_14_25 ();
 FILLCELL_X1 FILLER_14_27 ();
 FILLCELL_X2 FILLER_14_32 ();
 FILLCELL_X1 FILLER_14_41 ();
 FILLCELL_X1 FILLER_14_46 ();
 FILLCELL_X8 FILLER_14_87 ();
 FILLCELL_X4 FILLER_14_95 ();
 FILLCELL_X2 FILLER_14_99 ();
 FILLCELL_X1 FILLER_14_101 ();
 FILLCELL_X1 FILLER_14_106 ();
 FILLCELL_X1 FILLER_14_110 ();
 FILLCELL_X1 FILLER_14_118 ();
 FILLCELL_X4 FILLER_14_121 ();
 FILLCELL_X2 FILLER_14_125 ();
 FILLCELL_X8 FILLER_14_134 ();
 FILLCELL_X4 FILLER_14_142 ();
 FILLCELL_X4 FILLER_14_167 ();
 FILLCELL_X2 FILLER_14_171 ();
 FILLCELL_X1 FILLER_14_173 ();
 FILLCELL_X2 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_20 ();
 FILLCELL_X1 FILLER_15_22 ();
 FILLCELL_X1 FILLER_15_30 ();
 FILLCELL_X1 FILLER_15_35 ();
 FILLCELL_X1 FILLER_15_43 ();
 FILLCELL_X1 FILLER_15_52 ();
 FILLCELL_X1 FILLER_15_56 ();
 FILLCELL_X1 FILLER_15_68 ();
 FILLCELL_X1 FILLER_15_74 ();
 FILLCELL_X8 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_105 ();
 FILLCELL_X1 FILLER_15_109 ();
 FILLCELL_X1 FILLER_15_130 ();
 FILLCELL_X1 FILLER_15_135 ();
 FILLCELL_X4 FILLER_15_155 ();
 FILLCELL_X1 FILLER_15_159 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_13 ();
 FILLCELL_X8 FILLER_16_18 ();
 FILLCELL_X2 FILLER_16_26 ();
 FILLCELL_X1 FILLER_16_28 ();
 FILLCELL_X2 FILLER_16_46 ();
 FILLCELL_X1 FILLER_16_48 ();
 FILLCELL_X8 FILLER_16_57 ();
 FILLCELL_X4 FILLER_16_65 ();
 FILLCELL_X1 FILLER_16_69 ();
 FILLCELL_X16 FILLER_16_105 ();
 FILLCELL_X4 FILLER_16_121 ();
 FILLCELL_X2 FILLER_16_125 ();
 FILLCELL_X16 FILLER_16_131 ();
 FILLCELL_X4 FILLER_16_147 ();
 FILLCELL_X2 FILLER_16_151 ();
 FILLCELL_X8 FILLER_16_164 ();
 FILLCELL_X2 FILLER_16_172 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_5 ();
 FILLCELL_X1 FILLER_17_7 ();
 FILLCELL_X4 FILLER_17_11 ();
 FILLCELL_X4 FILLER_17_26 ();
 FILLCELL_X4 FILLER_17_34 ();
 FILLCELL_X2 FILLER_17_38 ();
 FILLCELL_X1 FILLER_17_40 ();
 FILLCELL_X8 FILLER_17_58 ();
 FILLCELL_X4 FILLER_17_83 ();
 FILLCELL_X2 FILLER_17_87 ();
 FILLCELL_X1 FILLER_17_89 ();
 FILLCELL_X8 FILLER_17_95 ();
 FILLCELL_X4 FILLER_17_103 ();
 FILLCELL_X2 FILLER_17_107 ();
 FILLCELL_X1 FILLER_17_109 ();
 FILLCELL_X8 FILLER_17_117 ();
 FILLCELL_X4 FILLER_17_125 ();
 FILLCELL_X2 FILLER_17_129 ();
 FILLCELL_X1 FILLER_17_131 ();
 FILLCELL_X4 FILLER_17_143 ();
 FILLCELL_X2 FILLER_17_147 ();
 FILLCELL_X4 FILLER_17_156 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_5 ();
 FILLCELL_X4 FILLER_18_28 ();
 FILLCELL_X2 FILLER_18_36 ();
 FILLCELL_X1 FILLER_18_38 ();
 FILLCELL_X8 FILLER_18_42 ();
 FILLCELL_X1 FILLER_18_50 ();
 FILLCELL_X8 FILLER_18_56 ();
 FILLCELL_X2 FILLER_18_64 ();
 FILLCELL_X4 FILLER_18_74 ();
 FILLCELL_X1 FILLER_18_78 ();
 FILLCELL_X8 FILLER_18_82 ();
 FILLCELL_X4 FILLER_18_90 ();
 FILLCELL_X2 FILLER_18_94 ();
 FILLCELL_X4 FILLER_18_117 ();
 FILLCELL_X4 FILLER_18_126 ();
 FILLCELL_X1 FILLER_18_130 ();
 FILLCELL_X4 FILLER_18_152 ();
 FILLCELL_X8 FILLER_18_160 ();
 FILLCELL_X4 FILLER_18_168 ();
 FILLCELL_X2 FILLER_18_172 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_9 ();
 FILLCELL_X4 FILLER_19_52 ();
 FILLCELL_X2 FILLER_19_56 ();
 FILLCELL_X1 FILLER_19_61 ();
 FILLCELL_X1 FILLER_19_84 ();
 FILLCELL_X1 FILLER_19_89 ();
 FILLCELL_X1 FILLER_19_97 ();
 FILLCELL_X8 FILLER_19_102 ();
 FILLCELL_X4 FILLER_19_110 ();
 FILLCELL_X16 FILLER_19_118 ();
 FILLCELL_X8 FILLER_19_134 ();
 FILLCELL_X4 FILLER_19_142 ();
 FILLCELL_X2 FILLER_19_146 ();
 FILLCELL_X1 FILLER_19_148 ();
 FILLCELL_X1 FILLER_19_153 ();
 FILLCELL_X2 FILLER_19_157 ();
 FILLCELL_X1 FILLER_19_159 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_17 ();
 FILLCELL_X1 FILLER_20_25 ();
 FILLCELL_X1 FILLER_20_29 ();
 FILLCELL_X8 FILLER_20_34 ();
 FILLCELL_X4 FILLER_20_42 ();
 FILLCELL_X4 FILLER_20_63 ();
 FILLCELL_X8 FILLER_20_69 ();
 FILLCELL_X4 FILLER_20_94 ();
 FILLCELL_X2 FILLER_20_98 ();
 FILLCELL_X1 FILLER_20_100 ();
 FILLCELL_X2 FILLER_20_105 ();
 FILLCELL_X2 FILLER_20_141 ();
 FILLCELL_X8 FILLER_20_167 ();
 FILLCELL_X2 FILLER_20_175 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X16 FILLER_21_32 ();
 FILLCELL_X4 FILLER_21_55 ();
 FILLCELL_X8 FILLER_21_66 ();
 FILLCELL_X8 FILLER_21_81 ();
 FILLCELL_X2 FILLER_21_96 ();
 FILLCELL_X2 FILLER_21_123 ();
 FILLCELL_X4 FILLER_21_142 ();
 FILLCELL_X16 FILLER_21_150 ();
 FILLCELL_X8 FILLER_21_166 ();
 FILLCELL_X2 FILLER_21_174 ();
 FILLCELL_X1 FILLER_21_176 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X2 FILLER_22_13 ();
 FILLCELL_X2 FILLER_22_32 ();
 FILLCELL_X1 FILLER_22_34 ();
 FILLCELL_X2 FILLER_22_56 ();
 FILLCELL_X1 FILLER_22_58 ();
 FILLCELL_X1 FILLER_22_63 ();
 FILLCELL_X1 FILLER_22_81 ();
 FILLCELL_X2 FILLER_22_86 ();
 FILLCELL_X4 FILLER_22_105 ();
 FILLCELL_X2 FILLER_22_109 ();
 FILLCELL_X1 FILLER_22_111 ();
 FILLCELL_X2 FILLER_22_136 ();
 FILLCELL_X8 FILLER_22_162 ();
 FILLCELL_X4 FILLER_22_170 ();
 FILLCELL_X2 FILLER_22_174 ();
 FILLCELL_X1 FILLER_22_176 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X8 FILLER_23_17 ();
 FILLCELL_X2 FILLER_23_25 ();
 FILLCELL_X1 FILLER_23_27 ();
 FILLCELL_X8 FILLER_23_35 ();
 FILLCELL_X4 FILLER_23_43 ();
 FILLCELL_X1 FILLER_23_47 ();
 FILLCELL_X2 FILLER_23_51 ();
 FILLCELL_X1 FILLER_23_53 ();
 FILLCELL_X2 FILLER_23_74 ();
 FILLCELL_X2 FILLER_23_79 ();
 FILLCELL_X4 FILLER_23_84 ();
 FILLCELL_X2 FILLER_23_92 ();
 FILLCELL_X2 FILLER_23_100 ();
 FILLCELL_X1 FILLER_23_102 ();
 FILLCELL_X8 FILLER_23_106 ();
 FILLCELL_X1 FILLER_23_114 ();
 FILLCELL_X8 FILLER_23_118 ();
 FILLCELL_X4 FILLER_23_126 ();
 FILLCELL_X2 FILLER_23_130 ();
 FILLCELL_X1 FILLER_23_132 ();
 FILLCELL_X8 FILLER_23_136 ();
 FILLCELL_X4 FILLER_23_144 ();
 FILLCELL_X2 FILLER_23_148 ();
 FILLCELL_X1 FILLER_23_150 ();
 FILLCELL_X16 FILLER_23_157 ();
 FILLCELL_X4 FILLER_23_173 ();
endmodule
