module non_restoring_divider (busy,
    clk,
    error,
    rst_n,
    start,
    valid,
    dividend,
    divisor,
    quotient,
    remainder);
 output busy;
 input clk;
 output error;
 input rst_n;
 input start;
 output valid;
 input [7:0] dividend;
 input [7:0] divisor;
 output [7:0] quotient;
 output [7:0] remainder;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire \div_reg[0] ;
 wire \div_reg[1] ;
 wire \div_reg[2] ;
 wire \div_reg[3] ;
 wire \div_reg[4] ;
 wire \div_reg[5] ;
 wire \div_reg[6] ;
 wire \div_reg[7] ;
 wire \iter[0] ;
 wire \iter[1] ;
 wire \iter[2] ;
 wire \iter[3] ;
 wire \quot[0] ;
 wire \quot[1] ;
 wire \quot[2] ;
 wire \quot[3] ;
 wire \quot[4] ;
 wire \quot[5] ;
 wire \quot[6] ;
 wire \quot[7] ;
 wire \rem[0] ;
 wire \rem[1] ;
 wire \rem[2] ;
 wire \rem[3] ;
 wire \rem[4] ;
 wire \rem[5] ;
 wire \rem[6] ;
 wire \rem[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net38;

 sky130_fd_sc_hd__clkbuf_2 _206_ (.A(\iter[2] ),
    .X(_049_));
 sky130_fd_sc_hd__nor2_1 _207_ (.A(\iter[0] ),
    .B(\iter[1] ),
    .Y(_050_));
 sky130_fd_sc_hd__nand2_1 _208_ (.A(\iter[3] ),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__mux4_1 _209_ (.A0(net5),
    .A1(net4),
    .A2(net3),
    .A3(net2),
    .S0(\iter[0] ),
    .S1(_159_),
    .X(_052_));
 sky130_fd_sc_hd__mux4_1 _210_ (.A0(net9),
    .A1(net8),
    .A2(net7),
    .A3(net6),
    .S0(\iter[0] ),
    .S1(_159_),
    .X(_053_));
 sky130_fd_sc_hd__mux2i_1 _211_ (.A0(_052_),
    .A1(_053_),
    .S(_160_),
    .Y(_054_));
 sky130_fd_sc_hd__nor3_1 _212_ (.A(_049_),
    .B(_160_),
    .C(_050_),
    .Y(_055_));
 sky130_fd_sc_hd__mux2_1 _213_ (.A0(_053_),
    .A1(_052_),
    .S(_160_),
    .X(_056_));
 sky130_fd_sc_hd__a22oi_1 _214_ (.A1(_052_),
    .A2(_055_),
    .B1(_056_),
    .B2(_049_),
    .Y(_057_));
 sky130_fd_sc_hd__o32a_1 _215_ (.A1(_049_),
    .A2(_051_),
    .A3(_054_),
    .B1(\iter[3] ),
    .B2(_057_),
    .X(_166_));
 sky130_fd_sc_hd__inv_1 _216_ (.A(_166_),
    .Y(_163_));
 sky130_fd_sc_hd__inv_1 _217_ (.A(\iter[0] ),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _218_ (.A(\div_reg[0] ),
    .Y(_162_));
 sky130_fd_sc_hd__inv_1 _219_ (.A(\div_reg[1] ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _220_ (.A(\div_reg[3] ),
    .Y(_173_));
 sky130_fd_sc_hd__inv_1 _221_ (.A(\div_reg[2] ),
    .Y(_179_));
 sky130_fd_sc_hd__inv_1 _222_ (.A(\div_reg[6] ),
    .Y(_188_));
 sky130_fd_sc_hd__inv_1 _223_ (.A(\div_reg[5] ),
    .Y(_194_));
 sky130_fd_sc_hd__inv_1 _224_ (.A(\div_reg[4] ),
    .Y(_200_));
 sky130_fd_sc_hd__inv_1 _225_ (.A(\iter[1] ),
    .Y(_157_));
 sky130_fd_sc_hd__inv_1 _226_ (.A(\rem[0] ),
    .Y(_152_));
 sky130_fd_sc_hd__inv_1 _227_ (.A(\rem[2] ),
    .Y(_176_));
 sky130_fd_sc_hd__inv_1 _228_ (.A(\rem[1] ),
    .Y(_182_));
 sky130_fd_sc_hd__inv_1 _229_ (.A(\rem[6] ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_1 _230_ (.A(\rem[5] ),
    .Y(_191_));
 sky130_fd_sc_hd__inv_1 _231_ (.A(\rem[4] ),
    .Y(_197_));
 sky130_fd_sc_hd__inv_1 _232_ (.A(\rem[3] ),
    .Y(_203_));
 sky130_fd_sc_hd__nor2_1 _233_ (.A(\state[1] ),
    .B(\state[0] ),
    .Y(_058_));
 sky130_fd_sc_hd__inv_1 _234_ (.A(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__nor2b_1 _235_ (.A(\state[1] ),
    .B_N(\state[0] ),
    .Y(_060_));
 sky130_fd_sc_hd__nor2b_1 _236_ (.A(_049_),
    .B_N(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__nand3b_4 _237_ (.A_N(\iter[3] ),
    .B(_158_),
    .C(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__clkbuf_4 _238_ (.A(_062_),
    .X(_063_));
 sky130_fd_sc_hd__nor4_2 _239_ (.A(net15),
    .B(net14),
    .C(net17),
    .D(net16),
    .Y(_064_));
 sky130_fd_sc_hd__nor4_2 _240_ (.A(net11),
    .B(net10),
    .C(net13),
    .D(net12),
    .Y(_065_));
 sky130_fd_sc_hd__nand2_1 _241_ (.A(net18),
    .B(_058_),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_4 _242_ (.A1(_064_),
    .A2(_065_),
    .B1(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net19),
    .A2(_059_),
    .A3(_063_),
    .B1(_067_),
    .X(_000_));
 sky130_fd_sc_hd__clkbuf_2 _244_ (.A(_067_),
    .X(_068_));
 sky130_fd_sc_hd__nand2_1 _245_ (.A(net10),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__o21ai_0 _246_ (.A1(_162_),
    .A2(_068_),
    .B1(_069_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _247_ (.A(net11),
    .B(_068_),
    .Y(_070_));
 sky130_fd_sc_hd__o21ai_0 _248_ (.A1(_168_),
    .A2(_068_),
    .B1(_070_),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(net12),
    .B(_068_),
    .Y(_071_));
 sky130_fd_sc_hd__o21ai_0 _250_ (.A1(_179_),
    .A2(_068_),
    .B1(_071_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _251_ (.A(net13),
    .B(_067_),
    .Y(_072_));
 sky130_fd_sc_hd__o21ai_0 _252_ (.A1(_173_),
    .A2(_068_),
    .B1(_072_),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _253_ (.A(net14),
    .B(_067_),
    .Y(_073_));
 sky130_fd_sc_hd__o21ai_0 _254_ (.A1(_200_),
    .A2(_068_),
    .B1(_073_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(net15),
    .B(_067_),
    .Y(_074_));
 sky130_fd_sc_hd__o21ai_0 _256_ (.A1(_194_),
    .A2(_068_),
    .B1(_074_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _257_ (.A(net16),
    .B(_067_),
    .Y(_075_));
 sky130_fd_sc_hd__o21ai_0 _258_ (.A1(_188_),
    .A2(_068_),
    .B1(_075_),
    .Y(_007_));
 sky130_fd_sc_hd__mux2_1 _259_ (.A0(\div_reg[7] ),
    .A1(net17),
    .S(_067_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(_064_),
    .B(_065_),
    .Y(_076_));
 sky130_fd_sc_hd__o2bb2ai_1 _261_ (.A1_N(net20),
    .A2_N(_059_),
    .B1(_066_),
    .B2(_076_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2b_1 _262_ (.A_N(\iter[3] ),
    .B(_158_),
    .Y(_077_));
 sky130_fd_sc_hd__o21ai_1 _263_ (.A1(_049_),
    .A2(_077_),
    .B1(_060_),
    .Y(_078_));
 sky130_fd_sc_hd__clkbuf_4 _264_ (.A(_078_),
    .X(_079_));
 sky130_fd_sc_hd__o21a_1 _265_ (.A1(_049_),
    .A2(_077_),
    .B1(_060_),
    .X(_080_));
 sky130_fd_sc_hd__buf_2 _266_ (.A(_080_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(_067_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__clkbuf_4 _268_ (.A(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nand2_1 _269_ (.A(\iter[0] ),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__o21ai_0 _270_ (.A1(\iter[0] ),
    .A2(_079_),
    .B1(_084_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _271_ (.A(_082_),
    .Y(_046_));
 sky130_fd_sc_hd__o22ai_1 _272_ (.A1(_159_),
    .A2(_079_),
    .B1(_046_),
    .B2(_157_),
    .Y(_011_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_160_),
    .B(_081_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _274_ (.A(_160_),
    .B(_079_),
    .Y(_086_));
 sky130_fd_sc_hd__o21ai_0 _275_ (.A1(_082_),
    .A2(_086_),
    .B1(_049_),
    .Y(_087_));
 sky130_fd_sc_hd__o21ai_0 _276_ (.A1(_049_),
    .A2(_085_),
    .B1(_087_),
    .Y(_012_));
 sky130_fd_sc_hd__nor2_1 _277_ (.A(_158_),
    .B(_050_),
    .Y(_088_));
 sky130_fd_sc_hd__o21ai_0 _278_ (.A1(_049_),
    .A2(_088_),
    .B1(_060_),
    .Y(_089_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(_046_),
    .A2(_089_),
    .B1(\iter[3] ),
    .Y(_090_));
 sky130_fd_sc_hd__a31oi_1 _280_ (.A1(\iter[3] ),
    .A2(_050_),
    .A3(_061_),
    .B1(_090_),
    .Y(_013_));
 sky130_fd_sc_hd__nand4_2 _281_ (.A(_187_),
    .B(_190_),
    .C(_196_),
    .D(_202_),
    .Y(_091_));
 sky130_fd_sc_hd__nand4_1 _282_ (.A(_170_),
    .B(_165_),
    .C(_175_),
    .D(_181_),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _283_ (.A(_187_),
    .B(_190_),
    .Y(_093_));
 sky130_fd_sc_hd__a21oi_1 _284_ (.A1(_204_),
    .A2(_196_),
    .B1(_198_),
    .Y(_094_));
 sky130_fd_sc_hd__a21oi_1 _285_ (.A1(_192_),
    .A2(_187_),
    .B1(_186_),
    .Y(_095_));
 sky130_fd_sc_hd__o21ai_2 _286_ (.A1(_093_),
    .A2(_094_),
    .B1(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2b_1 _287_ (.A(_164_),
    .B_N(_170_),
    .Y(_097_));
 sky130_fd_sc_hd__o211ai_1 _288_ (.A1(_171_),
    .A2(_097_),
    .B1(_175_),
    .C1(_181_),
    .Y(_098_));
 sky130_fd_sc_hd__a21oi_1 _289_ (.A1(_183_),
    .A2(_175_),
    .B1(_177_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _290_ (.A1(_098_),
    .A2(_099_),
    .B1(_091_),
    .Y(_100_));
 sky130_fd_sc_hd__o22ai_4 _291_ (.A1(_091_),
    .A2(_092_),
    .B1(_096_),
    .B2(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__nand2_1 _292_ (.A(_081_),
    .B(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__nand2_1 _293_ (.A(\quot[0] ),
    .B(_083_),
    .Y(_103_));
 sky130_fd_sc_hd__nand2_1 _294_ (.A(_102_),
    .B(_103_),
    .Y(_014_));
 sky130_fd_sc_hd__a22o_1 _295_ (.A1(\quot[0] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[1] ),
    .X(_015_));
 sky130_fd_sc_hd__a22o_1 _296_ (.A1(\quot[1] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[2] ),
    .X(_016_));
 sky130_fd_sc_hd__a22o_1 _297_ (.A1(\quot[2] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[3] ),
    .X(_017_));
 sky130_fd_sc_hd__a22o_1 _298_ (.A1(\quot[3] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[4] ),
    .X(_018_));
 sky130_fd_sc_hd__a22o_1 _299_ (.A1(\quot[4] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[5] ),
    .X(_019_));
 sky130_fd_sc_hd__a22o_1 _300_ (.A1(\quot[5] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[6] ),
    .X(_020_));
 sky130_fd_sc_hd__a22o_1 _301_ (.A1(\quot[6] ),
    .A2(_081_),
    .B1(_083_),
    .B2(\quot[7] ),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(\quot[0] ),
    .A1(net21),
    .S(_063_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\quot[1] ),
    .A1(net22),
    .S(_063_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _304_ (.A0(\quot[2] ),
    .A1(net23),
    .S(_063_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\quot[3] ),
    .A1(net24),
    .S(_062_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\quot[4] ),
    .A1(net25),
    .S(_062_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(\quot[5] ),
    .A1(net26),
    .S(_062_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\quot[6] ),
    .A1(net27),
    .S(_062_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\quot[7] ),
    .A1(net28),
    .S(_062_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(_166_),
    .A1(_165_),
    .S(_101_),
    .X(_104_));
 sky130_fd_sc_hd__o22ai_1 _311_ (.A1(_152_),
    .A2(_046_),
    .B1(_104_),
    .B2(_079_),
    .Y(_030_));
 sky130_fd_sc_hd__mux2i_1 _312_ (.A0(\rem[0] ),
    .A1(_155_),
    .S(_101_),
    .Y(_105_));
 sky130_fd_sc_hd__o22ai_1 _313_ (.A1(_182_),
    .A2(_046_),
    .B1(_105_),
    .B2(_079_),
    .Y(_031_));
 sky130_fd_sc_hd__xnor2_1 _314_ (.A(_154_),
    .B(_181_),
    .Y(_106_));
 sky130_fd_sc_hd__mux2i_1 _315_ (.A0(\rem[1] ),
    .A1(_106_),
    .S(_101_),
    .Y(_107_));
 sky130_fd_sc_hd__o22ai_1 _316_ (.A1(_176_),
    .A2(_046_),
    .B1(_107_),
    .B2(_079_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2b_1 _317_ (.A_N(_153_),
    .B(_170_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2b_1 _318_ (.A_N(_169_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__a211oi_1 _319_ (.A1(_181_),
    .A2(_109_),
    .B1(_180_),
    .C1(_175_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(_169_),
    .B(_180_),
    .Y(_111_));
 sky130_fd_sc_hd__o21ai_0 _321_ (.A1(_181_),
    .A2(_180_),
    .B1(_175_),
    .Y(_112_));
 sky130_fd_sc_hd__a21oi_1 _322_ (.A1(_108_),
    .A2(_111_),
    .B1(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__nor2_1 _323_ (.A(_110_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2i_1 _324_ (.A0(\rem[2] ),
    .A1(_114_),
    .S(_101_),
    .Y(_115_));
 sky130_fd_sc_hd__o22ai_1 _325_ (.A1(_203_),
    .A2(_046_),
    .B1(_115_),
    .B2(_079_),
    .Y(_033_));
 sky130_fd_sc_hd__o21ai_0 _326_ (.A1(_175_),
    .A2(_174_),
    .B1(_202_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2b_1 _327_ (.A(_154_),
    .B_N(_181_),
    .Y(_117_));
 sky130_fd_sc_hd__nor3_1 _328_ (.A(_174_),
    .B(_180_),
    .C(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__nor2_1 _329_ (.A(_202_),
    .B(_174_),
    .Y(_119_));
 sky130_fd_sc_hd__o21ai_0 _330_ (.A1(_180_),
    .A2(_117_),
    .B1(_175_),
    .Y(_120_));
 sky130_fd_sc_hd__a2bb2oi_1 _331_ (.A1_N(_116_),
    .A2_N(_118_),
    .B1(_119_),
    .B2(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__mux2i_1 _332_ (.A0(\rem[3] ),
    .A1(_121_),
    .S(_101_),
    .Y(_122_));
 sky130_fd_sc_hd__o22ai_1 _333_ (.A1(_197_),
    .A2(_046_),
    .B1(_122_),
    .B2(_079_),
    .Y(_034_));
 sky130_fd_sc_hd__o21ai_0 _334_ (.A1(_174_),
    .A2(_113_),
    .B1(_202_),
    .Y(_123_));
 sky130_fd_sc_hd__nand2b_1 _335_ (.A_N(_201_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__xnor2_1 _336_ (.A(_196_),
    .B(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o32ai_1 _337_ (.A1(_197_),
    .A2(_079_),
    .A3(_101_),
    .B1(_046_),
    .B2(_191_),
    .Y(_126_));
 sky130_fd_sc_hd__o21bai_1 _338_ (.A1(_102_),
    .A2(_125_),
    .B1_N(_126_),
    .Y(_035_));
 sky130_fd_sc_hd__o21bai_1 _339_ (.A1(_118_),
    .A2(_116_),
    .B1_N(_201_),
    .Y(_127_));
 sky130_fd_sc_hd__a21oi_1 _340_ (.A1(_196_),
    .A2(_127_),
    .B1(_195_),
    .Y(_128_));
 sky130_fd_sc_hd__xor2_1 _341_ (.A(_190_),
    .B(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o32ai_1 _342_ (.A1(_191_),
    .A2(_078_),
    .A3(_101_),
    .B1(_046_),
    .B2(_185_),
    .Y(_130_));
 sky130_fd_sc_hd__o21bai_1 _343_ (.A1(_102_),
    .A2(_129_),
    .B1_N(_130_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(\rem[6] ),
    .B(_101_),
    .Y(_131_));
 sky130_fd_sc_hd__a21oi_1 _345_ (.A1(_202_),
    .A2(_174_),
    .B1(_201_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2b_1 _346_ (.A(_132_),
    .B_N(_196_),
    .Y(_133_));
 sky130_fd_sc_hd__nand2_1 _347_ (.A(_196_),
    .B(_202_),
    .Y(_134_));
 sky130_fd_sc_hd__a211oi_1 _348_ (.A1(_108_),
    .A2(_111_),
    .B1(_112_),
    .C1(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__o31a_1 _349_ (.A1(_195_),
    .A2(_133_),
    .A3(_135_),
    .B1(_190_),
    .X(_136_));
 sky130_fd_sc_hd__o21ai_0 _350_ (.A1(_189_),
    .A2(_136_),
    .B1(_187_),
    .Y(_137_));
 sky130_fd_sc_hd__or3_1 _351_ (.A(_187_),
    .B(_189_),
    .C(_136_),
    .X(_138_));
 sky130_fd_sc_hd__a21boi_0 _352_ (.A1(_137_),
    .A2(_138_),
    .B1_N(_101_),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _353_ (.A(\rem[7] ),
    .B(_083_),
    .Y(_140_));
 sky130_fd_sc_hd__o31ai_1 _354_ (.A1(_079_),
    .A2(_131_),
    .A3(_139_),
    .B1(_140_),
    .Y(_037_));
 sky130_fd_sc_hd__buf_2 _355_ (.A(_062_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _356_ (.A(net29),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__o21ai_0 _357_ (.A1(_152_),
    .A2(_141_),
    .B1(_142_),
    .Y(_038_));
 sky130_fd_sc_hd__nand2_1 _358_ (.A(net30),
    .B(_063_),
    .Y(_143_));
 sky130_fd_sc_hd__o21ai_0 _359_ (.A1(_182_),
    .A2(_141_),
    .B1(_143_),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(net31),
    .B(_063_),
    .Y(_144_));
 sky130_fd_sc_hd__o21ai_0 _361_ (.A1(_176_),
    .A2(_141_),
    .B1(_144_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _362_ (.A(net32),
    .B(_063_),
    .Y(_145_));
 sky130_fd_sc_hd__o21ai_0 _363_ (.A1(_203_),
    .A2(_141_),
    .B1(_145_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(net33),
    .B(_063_),
    .Y(_146_));
 sky130_fd_sc_hd__o21ai_0 _365_ (.A1(_197_),
    .A2(_141_),
    .B1(_146_),
    .Y(_042_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(net34),
    .B(_063_),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_0 _367_ (.A1(_191_),
    .A2(_141_),
    .B1(_147_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _368_ (.A(net35),
    .B(_063_),
    .Y(_148_));
 sky130_fd_sc_hd__o21ai_0 _369_ (.A1(_185_),
    .A2(_141_),
    .B1(_148_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(\rem[7] ),
    .A1(net36),
    .S(_062_),
    .X(_045_));
 sky130_fd_sc_hd__nand2b_1 _371_ (.A_N(net18),
    .B(\state[1] ),
    .Y(_149_));
 sky130_fd_sc_hd__o21ai_0 _372_ (.A1(\state[0] ),
    .A2(_149_),
    .B1(_141_),
    .Y(_047_));
 sky130_fd_sc_hd__nand2b_1 _373_ (.A_N(\state[0] ),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__nand2_1 _374_ (.A(net37),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nand2_1 _375_ (.A(_141_),
    .B(_151_),
    .Y(_048_));
 sky130_fd_sc_hd__fa_1 _376_ (.A(\div_reg[1] ),
    .B(_152_),
    .CIN(_153_),
    .COUT(_154_),
    .SUM(_155_));
 sky130_fd_sc_hd__ha_1 _377_ (.A(_156_),
    .B(_157_),
    .COUT(_158_),
    .SUM(_159_));
 sky130_fd_sc_hd__ha_1 _378_ (.A(_156_),
    .B(_157_),
    .COUT(_160_),
    .SUM(_161_));
 sky130_fd_sc_hd__ha_1 _379_ (.A(_162_),
    .B(_163_),
    .COUT(_164_),
    .SUM(_165_));
 sky130_fd_sc_hd__ha_1 _380_ (.A(\div_reg[0] ),
    .B(_166_),
    .COUT(_153_),
    .SUM(_167_));
 sky130_fd_sc_hd__ha_1 _381_ (.A(_168_),
    .B(\rem[0] ),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__ha_1 _382_ (.A(\div_reg[1] ),
    .B(_152_),
    .COUT(_171_),
    .SUM(_172_));
 sky130_fd_sc_hd__ha_1 _383_ (.A(_173_),
    .B(\rem[2] ),
    .COUT(_174_),
    .SUM(_175_));
 sky130_fd_sc_hd__ha_1 _384_ (.A(\div_reg[3] ),
    .B(_176_),
    .COUT(_177_),
    .SUM(_178_));
 sky130_fd_sc_hd__ha_1 _385_ (.A(_179_),
    .B(\rem[1] ),
    .COUT(_180_),
    .SUM(_181_));
 sky130_fd_sc_hd__ha_1 _386_ (.A(\div_reg[2] ),
    .B(_182_),
    .COUT(_183_),
    .SUM(_184_));
 sky130_fd_sc_hd__ha_1 _387_ (.A(\div_reg[7] ),
    .B(_185_),
    .COUT(_186_),
    .SUM(_187_));
 sky130_fd_sc_hd__ha_1 _388_ (.A(_188_),
    .B(\rem[5] ),
    .COUT(_189_),
    .SUM(_190_));
 sky130_fd_sc_hd__ha_1 _389_ (.A(\div_reg[6] ),
    .B(_191_),
    .COUT(_192_),
    .SUM(_193_));
 sky130_fd_sc_hd__ha_2 _390_ (.A(_194_),
    .B(\rem[4] ),
    .COUT(_195_),
    .SUM(_196_));
 sky130_fd_sc_hd__ha_1 _391_ (.A(\div_reg[5] ),
    .B(_197_),
    .COUT(_198_),
    .SUM(_199_));
 sky130_fd_sc_hd__ha_1 _392_ (.A(_200_),
    .B(\rem[3] ),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__ha_1 _393_ (.A(\div_reg[4] ),
    .B(_203_),
    .COUT(_204_),
    .SUM(_205_));
 sky130_fd_sc_hd__dfrtp_1 \busy$_DFFE_PN0P_  (.D(_000_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[0]$_DFFE_PN0P_  (.D(_001_),
    .Q(\div_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[1]$_DFFE_PN0P_  (.D(_002_),
    .Q(\div_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[2]$_DFFE_PN0P_  (.D(_003_),
    .Q(\div_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[3]$_DFFE_PN0P_  (.D(_004_),
    .Q(\div_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[4]$_DFFE_PN0P_  (.D(_005_),
    .Q(\div_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[5]$_DFFE_PN0P_  (.D(_006_),
    .Q(\div_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[6]$_DFFE_PN0P_  (.D(_007_),
    .Q(\div_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \div_reg[7]$_DFFE_PN0P_  (.D(_008_),
    .Q(\div_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error$_DFFE_PN0P_  (.D(_009_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \iter[0]$_DFFE_PN0P_  (.D(_010_),
    .Q(\iter[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \iter[1]$_DFFE_PN0P_  (.D(_011_),
    .Q(\iter[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \iter[2]$_DFFE_PN0P_  (.D(_012_),
    .Q(\iter[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \iter[3]$_DFFE_PN0P_  (.D(_013_),
    .Q(\iter[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[0]$_DFFE_PN0P_  (.D(_014_),
    .Q(\quot[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[1]$_DFFE_PN0P_  (.D(_015_),
    .Q(\quot[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[2]$_DFFE_PN0P_  (.D(_016_),
    .Q(\quot[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[3]$_DFFE_PN0P_  (.D(_017_),
    .Q(\quot[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[4]$_DFFE_PN0P_  (.D(_018_),
    .Q(\quot[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[5]$_DFFE_PN0P_  (.D(_019_),
    .Q(\quot[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[6]$_DFFE_PN0P_  (.D(_020_),
    .Q(\quot[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quot[7]$_DFFE_PN0P_  (.D(_021_),
    .Q(\quot[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[0]$_DFFE_PN0P_  (.D(_022_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[2]$_DFFE_PN0P_  (.D(_024_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \quotient[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[0]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rem[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[1]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rem[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[2]$_DFFE_PN0P_  (.D(_032_),
    .Q(\rem[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[3]$_DFFE_PN0P_  (.D(_033_),
    .Q(\rem[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[4]$_DFFE_PN0P_  (.D(_034_),
    .Q(\rem[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[5]$_DFFE_PN0P_  (.D(_035_),
    .Q(\rem[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[6]$_DFFE_PN0P_  (.D(_036_),
    .Q(\rem[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rem[7]$_DFFE_PN0P_  (.D(_037_),
    .Q(\rem[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[0]$_DFFE_PN0P_  (.D(_038_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[1]$_DFFE_PN0P_  (.D(_039_),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[2]$_DFFE_PN0P_  (.D(_040_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[3]$_DFFE_PN0P_  (.D(_041_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[4]$_DFFE_PN0P_  (.D(_042_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[5]$_DFFE_PN0P_  (.D(_043_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[6]$_DFFE_PN0P_  (.D(_044_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \remainder[7]$_DFFE_PN0P_  (.D(_045_),
    .Q(net36),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_046_),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_047_),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid$_DFFE_PN0P_  (.D(_048_),
    .Q(net37),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net38),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_51 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(dividend[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dividend[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(dividend[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(dividend[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(dividend[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(dividend[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(dividend[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(dividend[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(divisor[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(divisor[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(divisor[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(divisor[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(divisor[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(divisor[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(divisor[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(divisor[7]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(start),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(busy));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(error));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(quotient[0]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(quotient[1]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(quotient[2]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(quotient[3]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(quotient[4]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(quotient[5]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(quotient[6]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(quotient[7]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(remainder[0]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(remainder[1]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(remainder[2]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(remainder[3]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(remainder[4]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(remainder[5]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(remainder[6]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(remainder[7]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net38));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
endmodule
