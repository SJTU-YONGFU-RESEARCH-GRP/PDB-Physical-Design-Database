module shift_register_right (clk,
    en,
    load,
    rst_n,
    serial_in,
    serial_out,
    parallel_in,
    parallel_out);
 input clk;
 input en;
 input load;
 input rst_n;
 input serial_in;
 output serial_out;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X2 _35_ (.A(rst_n),
    .Z(_08_));
 BUF_X4 _36_ (.A(en),
    .Z(_09_));
 MUX2_X1 _37_ (.A(net18),
    .B(net11),
    .S(_09_),
    .Z(_10_));
 CLKBUF_X3 _38_ (.A(load),
    .Z(_11_));
 MUX2_X1 _39_ (.A(_10_),
    .B(net1),
    .S(_11_),
    .Z(_12_));
 AND2_X1 _40_ (.A1(_08_),
    .A2(_12_),
    .ZN(_00_));
 MUX2_X1 _41_ (.A(net11),
    .B(net12),
    .S(_09_),
    .Z(_13_));
 MUX2_X1 _42_ (.A(_13_),
    .B(net2),
    .S(_11_),
    .Z(_14_));
 AND2_X1 _43_ (.A1(_08_),
    .A2(_14_),
    .ZN(_01_));
 MUX2_X1 _44_ (.A(net12),
    .B(net13),
    .S(_09_),
    .Z(_15_));
 MUX2_X1 _45_ (.A(_15_),
    .B(net3),
    .S(_11_),
    .Z(_16_));
 AND2_X1 _46_ (.A1(_08_),
    .A2(_16_),
    .ZN(_02_));
 MUX2_X1 _47_ (.A(net13),
    .B(net14),
    .S(_09_),
    .Z(_17_));
 MUX2_X1 _48_ (.A(_17_),
    .B(net4),
    .S(_11_),
    .Z(_18_));
 AND2_X1 _49_ (.A1(_08_),
    .A2(_18_),
    .ZN(_03_));
 MUX2_X1 _50_ (.A(net14),
    .B(net15),
    .S(_09_),
    .Z(_19_));
 MUX2_X1 _51_ (.A(_19_),
    .B(net5),
    .S(_11_),
    .Z(_20_));
 AND2_X1 _52_ (.A1(_08_),
    .A2(_20_),
    .ZN(_04_));
 MUX2_X1 _53_ (.A(net15),
    .B(net16),
    .S(_09_),
    .Z(_21_));
 MUX2_X1 _54_ (.A(_21_),
    .B(net6),
    .S(_11_),
    .Z(_22_));
 AND2_X1 _55_ (.A1(_08_),
    .A2(_22_),
    .ZN(_05_));
 MUX2_X1 _56_ (.A(net16),
    .B(net17),
    .S(_09_),
    .Z(_23_));
 MUX2_X1 _57_ (.A(_23_),
    .B(net7),
    .S(_11_),
    .Z(_24_));
 AND2_X1 _58_ (.A1(_08_),
    .A2(_24_),
    .ZN(_06_));
 MUX2_X1 _59_ (.A(net17),
    .B(net9),
    .S(_09_),
    .Z(_25_));
 MUX2_X1 _60_ (.A(_25_),
    .B(net8),
    .S(_11_),
    .Z(_26_));
 AND2_X1 _61_ (.A1(_08_),
    .A2(_26_),
    .ZN(_07_));
 BUF_X1 _62_ (.A(net18),
    .Z(net10));
 DFF_X1 \parallel_out[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_34_));
 DFF_X1 \parallel_out[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_33_));
 DFF_X1 \parallel_out[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net12),
    .QN(_32_));
 DFF_X1 \parallel_out[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_31_));
 DFF_X1 \parallel_out[4]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_30_));
 DFF_X1 \parallel_out[5]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net15),
    .QN(_29_));
 DFF_X1 \parallel_out[6]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_28_));
 DFF_X1 \parallel_out[7]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_27_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_57 ();
 BUF_X1 input1 (.A(parallel_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(parallel_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(parallel_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(parallel_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(parallel_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(parallel_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(parallel_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(parallel_in[7]),
    .Z(net8));
 BUF_X1 input9 (.A(serial_in),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(parallel_out[0]));
 BUF_X1 output11 (.A(net11),
    .Z(parallel_out[1]));
 BUF_X1 output12 (.A(net12),
    .Z(parallel_out[2]));
 BUF_X1 output13 (.A(net13),
    .Z(parallel_out[3]));
 BUF_X1 output14 (.A(net14),
    .Z(parallel_out[4]));
 BUF_X1 output15 (.A(net15),
    .Z(parallel_out[5]));
 BUF_X1 output16 (.A(net16),
    .Z(parallel_out[6]));
 BUF_X1 output17 (.A(net17),
    .Z(parallel_out[7]));
 BUF_X1 output18 (.A(net18),
    .Z(serial_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X32 FILLER_0_92 ();
 FILLCELL_X32 FILLER_0_124 ();
 FILLCELL_X32 FILLER_0_156 ();
 FILLCELL_X16 FILLER_0_188 ();
 FILLCELL_X8 FILLER_0_204 ();
 FILLCELL_X2 FILLER_0_212 ();
 FILLCELL_X1 FILLER_0_214 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X16 FILLER_1_193 ();
 FILLCELL_X4 FILLER_1_209 ();
 FILLCELL_X2 FILLER_1_213 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X16 FILLER_2_193 ();
 FILLCELL_X4 FILLER_2_209 ();
 FILLCELL_X2 FILLER_2_213 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X16 FILLER_3_193 ();
 FILLCELL_X4 FILLER_3_209 ();
 FILLCELL_X2 FILLER_3_213 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X16 FILLER_4_193 ();
 FILLCELL_X4 FILLER_4_209 ();
 FILLCELL_X2 FILLER_4_213 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X16 FILLER_5_193 ();
 FILLCELL_X4 FILLER_5_209 ();
 FILLCELL_X2 FILLER_5_213 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X16 FILLER_6_193 ();
 FILLCELL_X4 FILLER_6_209 ();
 FILLCELL_X2 FILLER_6_213 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X16 FILLER_7_193 ();
 FILLCELL_X4 FILLER_7_209 ();
 FILLCELL_X2 FILLER_7_213 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X16 FILLER_8_193 ();
 FILLCELL_X4 FILLER_8_209 ();
 FILLCELL_X2 FILLER_8_213 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X16 FILLER_9_193 ();
 FILLCELL_X4 FILLER_9_209 ();
 FILLCELL_X2 FILLER_9_213 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X16 FILLER_10_193 ();
 FILLCELL_X4 FILLER_10_209 ();
 FILLCELL_X2 FILLER_10_213 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_161 ();
 FILLCELL_X2 FILLER_11_177 ();
 FILLCELL_X16 FILLER_11_196 ();
 FILLCELL_X2 FILLER_11_212 ();
 FILLCELL_X1 FILLER_11_214 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_5 ();
 FILLCELL_X1 FILLER_12_7 ();
 FILLCELL_X16 FILLER_12_49 ();
 FILLCELL_X2 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_102 ();
 FILLCELL_X32 FILLER_12_134 ();
 FILLCELL_X4 FILLER_12_166 ();
 FILLCELL_X2 FILLER_12_170 ();
 FILLCELL_X2 FILLER_12_187 ();
 FILLCELL_X4 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_5 ();
 FILLCELL_X32 FILLER_13_11 ();
 FILLCELL_X32 FILLER_13_43 ();
 FILLCELL_X32 FILLER_13_75 ();
 FILLCELL_X32 FILLER_13_107 ();
 FILLCELL_X16 FILLER_13_139 ();
 FILLCELL_X8 FILLER_13_155 ();
 FILLCELL_X1 FILLER_13_163 ();
 FILLCELL_X4 FILLER_13_188 ();
 FILLCELL_X1 FILLER_13_192 ();
 FILLCELL_X8 FILLER_13_200 ();
 FILLCELL_X4 FILLER_13_208 ();
 FILLCELL_X2 FILLER_13_212 ();
 FILLCELL_X1 FILLER_13_214 ();
 FILLCELL_X8 FILLER_14_11 ();
 FILLCELL_X2 FILLER_14_19 ();
 FILLCELL_X2 FILLER_14_28 ();
 FILLCELL_X1 FILLER_14_30 ();
 FILLCELL_X16 FILLER_14_48 ();
 FILLCELL_X8 FILLER_14_64 ();
 FILLCELL_X16 FILLER_14_77 ();
 FILLCELL_X8 FILLER_14_93 ();
 FILLCELL_X4 FILLER_14_101 ();
 FILLCELL_X2 FILLER_14_105 ();
 FILLCELL_X1 FILLER_14_107 ();
 FILLCELL_X16 FILLER_14_113 ();
 FILLCELL_X8 FILLER_14_129 ();
 FILLCELL_X4 FILLER_14_137 ();
 FILLCELL_X2 FILLER_14_141 ();
 FILLCELL_X16 FILLER_14_148 ();
 FILLCELL_X8 FILLER_14_164 ();
 FILLCELL_X4 FILLER_14_172 ();
 FILLCELL_X2 FILLER_14_176 ();
 FILLCELL_X1 FILLER_14_178 ();
 FILLCELL_X8 FILLER_14_183 ();
 FILLCELL_X2 FILLER_14_191 ();
 FILLCELL_X1 FILLER_14_193 ();
 FILLCELL_X4 FILLER_14_206 ();
 FILLCELL_X2 FILLER_14_210 ();
 FILLCELL_X2 FILLER_15_7 ();
 FILLCELL_X32 FILLER_15_37 ();
 FILLCELL_X32 FILLER_15_69 ();
 FILLCELL_X32 FILLER_15_101 ();
 FILLCELL_X32 FILLER_15_133 ();
 FILLCELL_X8 FILLER_15_165 ();
 FILLCELL_X2 FILLER_15_173 ();
 FILLCELL_X1 FILLER_15_175 ();
 FILLCELL_X4 FILLER_15_200 ();
 FILLCELL_X2 FILLER_15_204 ();
 FILLCELL_X2 FILLER_15_212 ();
 FILLCELL_X1 FILLER_15_214 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_5 ();
 FILLCELL_X1 FILLER_16_7 ();
 FILLCELL_X2 FILLER_16_14 ();
 FILLCELL_X1 FILLER_16_16 ();
 FILLCELL_X1 FILLER_16_28 ();
 FILLCELL_X32 FILLER_16_36 ();
 FILLCELL_X32 FILLER_16_68 ();
 FILLCELL_X32 FILLER_16_100 ();
 FILLCELL_X32 FILLER_16_132 ();
 FILLCELL_X8 FILLER_16_164 ();
 FILLCELL_X4 FILLER_16_172 ();
 FILLCELL_X2 FILLER_16_176 ();
 FILLCELL_X1 FILLER_16_206 ();
 FILLCELL_X2 FILLER_16_210 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X16 FILLER_17_193 ();
 FILLCELL_X2 FILLER_17_212 ();
 FILLCELL_X1 FILLER_17_214 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X16 FILLER_18_193 ();
 FILLCELL_X4 FILLER_18_209 ();
 FILLCELL_X2 FILLER_18_213 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X16 FILLER_19_193 ();
 FILLCELL_X4 FILLER_19_209 ();
 FILLCELL_X2 FILLER_19_213 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X16 FILLER_20_193 ();
 FILLCELL_X4 FILLER_20_209 ();
 FILLCELL_X2 FILLER_20_213 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X16 FILLER_21_193 ();
 FILLCELL_X4 FILLER_21_209 ();
 FILLCELL_X2 FILLER_21_213 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X16 FILLER_22_193 ();
 FILLCELL_X4 FILLER_22_209 ();
 FILLCELL_X2 FILLER_22_213 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X16 FILLER_23_193 ();
 FILLCELL_X4 FILLER_23_209 ();
 FILLCELL_X2 FILLER_23_213 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X16 FILLER_24_193 ();
 FILLCELL_X4 FILLER_24_209 ();
 FILLCELL_X2 FILLER_24_213 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X4 FILLER_25_209 ();
 FILLCELL_X2 FILLER_25_213 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X16 FILLER_26_193 ();
 FILLCELL_X4 FILLER_26_209 ();
 FILLCELL_X2 FILLER_26_213 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X16 FILLER_27_193 ();
 FILLCELL_X4 FILLER_27_209 ();
 FILLCELL_X2 FILLER_27_213 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X16 FILLER_28_193 ();
 FILLCELL_X4 FILLER_28_209 ();
 FILLCELL_X2 FILLER_28_213 ();
endmodule
