module ddr_controller (clk,
    cmd_ready,
    cmd_valid,
    cmd_write,
    init_done,
    phy_cas_n,
    phy_cke,
    phy_clk,
    phy_cs_n,
    phy_odt,
    phy_ras_n,
    phy_reset_n,
    phy_we_n,
    rd_ready,
    rd_valid,
    rst_n,
    wr_ready,
    wr_valid,
    cmd_addr,
    cmd_burst_len,
    phy_addr,
    phy_bank,
    phy_bank_group,
    phy_dm,
    phy_dq,
    phy_dqs_n,
    phy_dqs_p,
    rd_data,
    state,
    wr_data,
    wr_mask);
 input clk;
 output cmd_ready;
 input cmd_valid;
 input cmd_write;
 output init_done;
 output phy_cas_n;
 output phy_cke;
 input phy_clk;
 output phy_cs_n;
 output phy_odt;
 output phy_ras_n;
 output phy_reset_n;
 output phy_we_n;
 input rd_ready;
 output rd_valid;
 input rst_n;
 output wr_ready;
 input wr_valid;
 input [27:0] cmd_addr;
 input [3:0] cmd_burst_len;
 output [13:0] phy_addr;
 output [2:0] phy_bank;
 output [1:0] phy_bank_group;
 output [7:0] phy_dm;
 inout [63:0] phy_dq;
 inout [7:0] phy_dqs_n;
 inout [7:0] phy_dqs_p;
 output [63:0] rd_data;
 output [1:0] state;
 input [63:0] wr_data;
 input [7:0] wr_mask;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire clknet_0_clk;
 wire net212;
 wire _0670_;
 wire \active_row[0][0] ;
 wire \active_row[0][10] ;
 wire \active_row[0][11] ;
 wire \active_row[0][12] ;
 wire \active_row[0][13] ;
 wire \active_row[0][1] ;
 wire \active_row[0][2] ;
 wire \active_row[0][3] ;
 wire \active_row[0][4] ;
 wire \active_row[0][5] ;
 wire \active_row[0][6] ;
 wire \active_row[0][7] ;
 wire \active_row[0][8] ;
 wire \active_row[0][9] ;
 wire \active_row[1][0] ;
 wire \active_row[1][10] ;
 wire \active_row[1][11] ;
 wire \active_row[1][12] ;
 wire \active_row[1][13] ;
 wire \active_row[1][1] ;
 wire \active_row[1][2] ;
 wire \active_row[1][3] ;
 wire \active_row[1][4] ;
 wire \active_row[1][5] ;
 wire \active_row[1][6] ;
 wire \active_row[1][7] ;
 wire \active_row[1][8] ;
 wire \active_row[1][9] ;
 wire \active_row[2][0] ;
 wire \active_row[2][10] ;
 wire \active_row[2][11] ;
 wire \active_row[2][12] ;
 wire \active_row[2][13] ;
 wire \active_row[2][1] ;
 wire \active_row[2][2] ;
 wire \active_row[2][3] ;
 wire \active_row[2][4] ;
 wire \active_row[2][5] ;
 wire \active_row[2][6] ;
 wire \active_row[2][7] ;
 wire \active_row[2][8] ;
 wire \active_row[2][9] ;
 wire \active_row[3][0] ;
 wire \active_row[3][10] ;
 wire \active_row[3][11] ;
 wire \active_row[3][12] ;
 wire \active_row[3][13] ;
 wire \active_row[3][1] ;
 wire \active_row[3][2] ;
 wire \active_row[3][3] ;
 wire \active_row[3][4] ;
 wire \active_row[3][5] ;
 wire \active_row[3][6] ;
 wire \active_row[3][7] ;
 wire \active_row[3][8] ;
 wire \active_row[3][9] ;
 wire \active_row[4][0] ;
 wire \active_row[4][10] ;
 wire \active_row[4][11] ;
 wire \active_row[4][12] ;
 wire \active_row[4][13] ;
 wire \active_row[4][1] ;
 wire \active_row[4][2] ;
 wire \active_row[4][3] ;
 wire \active_row[4][4] ;
 wire \active_row[4][5] ;
 wire \active_row[4][6] ;
 wire \active_row[4][7] ;
 wire \active_row[4][8] ;
 wire \active_row[4][9] ;
 wire \active_row[5][0] ;
 wire \active_row[5][10] ;
 wire \active_row[5][11] ;
 wire \active_row[5][12] ;
 wire \active_row[5][13] ;
 wire \active_row[5][1] ;
 wire \active_row[5][2] ;
 wire \active_row[5][3] ;
 wire \active_row[5][4] ;
 wire \active_row[5][5] ;
 wire \active_row[5][6] ;
 wire \active_row[5][7] ;
 wire \active_row[5][8] ;
 wire \active_row[5][9] ;
 wire \active_row[6][0] ;
 wire \active_row[6][10] ;
 wire \active_row[6][11] ;
 wire \active_row[6][12] ;
 wire \active_row[6][13] ;
 wire \active_row[6][1] ;
 wire \active_row[6][2] ;
 wire \active_row[6][3] ;
 wire \active_row[6][4] ;
 wire \active_row[6][5] ;
 wire \active_row[6][6] ;
 wire \active_row[6][7] ;
 wire \active_row[6][8] ;
 wire \active_row[6][9] ;
 wire \active_row[7][0] ;
 wire \active_row[7][10] ;
 wire \active_row[7][11] ;
 wire \active_row[7][12] ;
 wire \active_row[7][13] ;
 wire \active_row[7][1] ;
 wire \active_row[7][2] ;
 wire \active_row[7][3] ;
 wire \active_row[7][4] ;
 wire \active_row[7][5] ;
 wire \active_row[7][6] ;
 wire \active_row[7][7] ;
 wire \active_row[7][8] ;
 wire \active_row[7][9] ;
 wire \bank_active[0] ;
 wire \bank_active[1] ;
 wire \bank_active[2] ;
 wire \bank_active[3] ;
 wire \bank_active[4] ;
 wire \bank_active[5] ;
 wire \bank_active[6] ;
 wire \bank_active[7] ;
 wire \burst_counter[0] ;
 wire \burst_counter[1] ;
 wire \burst_counter[2] ;
 wire \burst_counter[3] ;
 wire cmd_reg_valid;
 wire \init_state[0] ;
 wire \init_state[1] ;
 wire \init_state[2] ;
 wire \init_state[3] ;
 wire \init_state[4] ;
 wire \init_state[5] ;
 wire \init_state[6] ;
 wire \init_state[7] ;
 wire \refresh_counter[0] ;
 wire \refresh_counter[10] ;
 wire \refresh_counter[11] ;
 wire \refresh_counter[12] ;
 wire \refresh_counter[13] ;
 wire \refresh_counter[14] ;
 wire \refresh_counter[15] ;
 wire \refresh_counter[1] ;
 wire \refresh_counter[2] ;
 wire \refresh_counter[3] ;
 wire \refresh_counter[4] ;
 wire \refresh_counter[5] ;
 wire \refresh_counter[6] ;
 wire \refresh_counter[7] ;
 wire \refresh_counter[8] ;
 wire \refresh_counter[9] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[1] ;
 wire \timer[2] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net223;

 sky130_fd_sc_hd__buf_2 _0671_ (.A(_0660_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _0672_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_0051_));
 sky130_fd_sc_hd__nor2_2 _0673_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .Y(_0052_));
 sky130_fd_sc_hd__and3_1 _0674_ (.A(_0654_),
    .B(_0051_),
    .C(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__or4_2 _0675_ (.A(\timer[7] ),
    .B(\timer[9] ),
    .C(\timer[8] ),
    .D(\timer[10] ),
    .X(_0054_));
 sky130_fd_sc_hd__or2_1 _0676_ (.A(\timer[6] ),
    .B(\timer[11] ),
    .X(_0055_));
 sky130_fd_sc_hd__or4_2 _0677_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[14] ),
    .D(\timer[15] ),
    .X(_0056_));
 sky130_fd_sc_hd__nor3_2 _0678_ (.A(_0054_),
    .B(_0055_),
    .C(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__and3_1 _0679_ (.A(_0050_),
    .B(_0053_),
    .C(_0057_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_2 _0680_ (.A(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(\init_state[4] ),
    .B(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__clkbuf_4 _0682_ (.A(_0050_),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_4 _0683_ (.A(_0061_),
    .X(_0062_));
 sky130_fd_sc_hd__nand3_4 _0684_ (.A(_0654_),
    .B(_0051_),
    .C(_0052_),
    .Y(_0063_));
 sky130_fd_sc_hd__or3_2 _0685_ (.A(_0054_),
    .B(_0055_),
    .C(_0056_),
    .X(_0064_));
 sky130_fd_sc_hd__nor2_1 _0686_ (.A(_0063_),
    .B(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__clkbuf_4 _0687_ (.A(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_4 _0688_ (.A(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_2 _0689_ (.A(_0062_),
    .B(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _0690_ (.A(\init_state[2] ),
    .B(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_1 _0691_ (.A(_0060_),
    .B(_0069_),
    .Y(_0003_));
 sky130_fd_sc_hd__clkbuf_4 _0692_ (.A(_0662_),
    .X(_0070_));
 sky130_fd_sc_hd__and3_2 _0693_ (.A(net36),
    .B(_0070_),
    .C(_0067_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_4 _0694_ (.A(_0631_),
    .B(_0071_),
    .X(_0012_));
 sky130_fd_sc_hd__inv_1 _0695_ (.A(net120),
    .Y(_0628_));
 sky130_fd_sc_hd__and3_4 _0696_ (.A(_0628_),
    .B(_0626_),
    .C(_0071_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _0697_ (.A(\init_state[5] ),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _0698_ (.A(_0072_),
    .B(_0059_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(\init_state[3] ),
    .B(_0068_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _0700_ (.A(_0073_),
    .B(_0074_),
    .Y(_0004_));
 sky130_fd_sc_hd__and3_4 _0701_ (.A(_0628_),
    .B(_0622_),
    .C(_0071_),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(\init_state[0] ),
    .B(_0059_),
    .Y(_0075_));
 sky130_fd_sc_hd__nand2_1 _0703_ (.A(\init_state[4] ),
    .B(_0068_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand2_1 _0704_ (.A(_0075_),
    .B(_0076_),
    .Y(_0005_));
 sky130_fd_sc_hd__and3_4 _0705_ (.A(_0628_),
    .B(_0624_),
    .C(_0071_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_4 _0706_ (.A(_0629_),
    .B(_0071_),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_1 _0707_ (.A(\init_state[1] ),
    .B(_0059_),
    .Y(_0077_));
 sky130_fd_sc_hd__nand2_1 _0708_ (.A(_0072_),
    .B(_0068_),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_1 _0709_ (.A(_0077_),
    .B(_0078_),
    .Y(_0006_));
 sky130_fd_sc_hd__and3_4 _0710_ (.A(net120),
    .B(_0624_),
    .C(_0071_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2b_1 _0711_ (.A(_0059_),
    .B_N(\init_state[0] ),
    .Y(_0001_));
 sky130_fd_sc_hd__and3_4 _0712_ (.A(net120),
    .B(_0626_),
    .C(_0071_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _0713_ (.A(\init_state[6] ),
    .B(_0059_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _0714_ (.A(\init_state[1] ),
    .B(_0068_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(_0079_),
    .B(_0080_),
    .Y(_0002_));
 sky130_fd_sc_hd__and3_4 _0716_ (.A(net120),
    .B(_0622_),
    .C(_0071_),
    .X(_0010_));
 sky130_fd_sc_hd__nand2_1 _0717_ (.A(\init_state[2] ),
    .B(_0059_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _0718_ (.A(\init_state[6] ),
    .B(_0068_),
    .Y(_0082_));
 sky130_fd_sc_hd__nand2_1 _0719_ (.A(_0081_),
    .B(_0082_),
    .Y(_0007_));
 sky130_fd_sc_hd__a21o_1 _0720_ (.A1(\init_state[3] ),
    .A2(_0059_),
    .B1(\init_state[7] ),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _0721_ (.A(_0666_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _0722_ (.A(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_4 _0723_ (.A(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2b_1 _0724_ (.A(net121),
    .B_N(net131),
    .Y(_0086_));
 sky130_fd_sc_hd__and3_4 _0725_ (.A(_0085_),
    .B(net133),
    .C(_0086_),
    .X(_0017_));
 sky130_fd_sc_hd__inv_1 _0726_ (.A(\burst_counter[0] ),
    .Y(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _0727_ (.A(net4),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_4 _0728_ (.A(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__buf_6 _0729_ (.A(cmd_addr[12]),
    .X(_0089_));
 sky130_fd_sc_hd__buf_6 _0730_ (.A(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__buf_6 _0731_ (.A(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__buf_6 _0732_ (.A(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__buf_4 _0733_ (.A(net3),
    .X(_0093_));
 sky130_fd_sc_hd__buf_6 _0734_ (.A(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__nor3b_1 _0735_ (.A(_0088_),
    .B(_0092_),
    .C_N(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_2 _0736_ (.A(_0088_),
    .B(_0092_),
    .Y(_0096_));
 sky130_fd_sc_hd__buf_6 _0737_ (.A(_0093_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2i_1 _0738_ (.A0(\active_row[6][9] ),
    .A1(\active_row[7][9] ),
    .S(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__o2bb2ai_1 _0739_ (.A1_N(\active_row[1][9] ),
    .A2_N(_0095_),
    .B1(_0096_),
    .B2(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_1 _0740_ (.A(_0089_),
    .Y(_0100_));
 sky130_fd_sc_hd__buf_4 _0741_ (.A(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__nor2b_1 _0742_ (.A(_0091_),
    .B_N(\active_row[4][9] ),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_1 _0743_ (.A(net4),
    .Y(_0103_));
 sky130_fd_sc_hd__buf_4 _0744_ (.A(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__clkinv_4 _0745_ (.A(_0093_),
    .Y(_0105_));
 sky130_fd_sc_hd__o221a_1 _0746_ (.A1(_0101_),
    .A2(\active_row[2][9] ),
    .B1(_0102_),
    .B2(_0104_),
    .C1(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_6 _0747_ (.A(_0091_),
    .X(_0107_));
 sky130_fd_sc_hd__inv_1 _0748_ (.A(\active_row[5][9] ),
    .Y(_0108_));
 sky130_fd_sc_hd__nand2_4 _0749_ (.A(_0088_),
    .B(_0097_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_1 _0750_ (.A(_0107_),
    .B(\active_row[3][9] ),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2b_4 _0751_ (.A_N(net4),
    .B(net3),
    .Y(_0111_));
 sky130_fd_sc_hd__o32ai_4 _0752_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0109_),
    .B1(_0110_),
    .B2(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__or3_1 _0753_ (.A(_0087_),
    .B(_0093_),
    .C(_0090_),
    .X(_0113_));
 sky130_fd_sc_hd__buf_4 _0754_ (.A(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__o32ai_4 _0755_ (.A1(_0099_),
    .A2(_0106_),
    .A3(_0112_),
    .B1(_0114_),
    .B2(\active_row[0][9] ),
    .Y(_0115_));
 sky130_fd_sc_hd__xor2_1 _0756_ (.A(net15),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2i_1 _0757_ (.A0(\active_row[6][3] ),
    .A1(\active_row[7][3] ),
    .S(_0097_),
    .Y(_0117_));
 sky130_fd_sc_hd__o2bb2ai_1 _0758_ (.A1_N(\active_row[1][3] ),
    .A2_N(_0095_),
    .B1(_0096_),
    .B2(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2b_1 _0759_ (.A(_0091_),
    .B_N(\active_row[4][3] ),
    .Y(_0119_));
 sky130_fd_sc_hd__o221a_1 _0760_ (.A1(_0101_),
    .A2(\active_row[2][3] ),
    .B1(_0119_),
    .B2(_0104_),
    .C1(_0105_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_6 _0761_ (.A(_0092_),
    .X(_0121_));
 sky130_fd_sc_hd__inv_1 _0762_ (.A(\active_row[5][3] ),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_1 _0763_ (.A(_0121_),
    .B(\active_row[3][3] ),
    .Y(_0123_));
 sky130_fd_sc_hd__o32ai_4 _0764_ (.A1(_0121_),
    .A2(_0122_),
    .A3(_0109_),
    .B1(_0123_),
    .B2(_0111_),
    .Y(_0124_));
 sky130_fd_sc_hd__o32ai_4 _0765_ (.A1(_0118_),
    .A2(_0120_),
    .A3(_0124_),
    .B1(_0114_),
    .B2(\active_row[0][3] ),
    .Y(_0125_));
 sky130_fd_sc_hd__xor2_1 _0766_ (.A(net8),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_1 _0767_ (.A(_0116_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__mux2i_1 _0768_ (.A0(\active_row[1][2] ),
    .A1(\active_row[3][2] ),
    .S(_0090_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand3b_1 _0769_ (.A_N(_0090_),
    .B(\active_row[5][2] ),
    .C(_0087_),
    .Y(_0129_));
 sky130_fd_sc_hd__o21ai_0 _0770_ (.A1(_0087_),
    .A2(_0128_),
    .B1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__and2_0 _0771_ (.A(net4),
    .B(_0089_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(\active_row[6][2] ),
    .A1(\active_row[7][2] ),
    .S(net3),
    .X(_0132_));
 sky130_fd_sc_hd__nand2b_1 _0773_ (.A_N(\active_row[2][2] ),
    .B(_0089_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_2 _0774_ (.A(net4),
    .B(net3),
    .Y(_0134_));
 sky130_fd_sc_hd__nor2_1 _0775_ (.A(_0093_),
    .B(_0090_),
    .Y(_0135_));
 sky130_fd_sc_hd__a222oi_1 _0776_ (.A1(_0131_),
    .A2(_0132_),
    .B1(_0133_),
    .B2(_0134_),
    .C1(_0135_),
    .C2(\active_row[4][2] ),
    .Y(_0136_));
 sky130_fd_sc_hd__a21boi_2 _0777_ (.A1(_0094_),
    .A2(_0130_),
    .B1_N(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__nor2_1 _0778_ (.A(\active_row[0][2] ),
    .B(_0113_),
    .Y(_0138_));
 sky130_fd_sc_hd__or3_1 _0779_ (.A(net7),
    .B(_0137_),
    .C(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _0780_ (.A(net7),
    .B(_0137_),
    .Y(_0140_));
 sky130_fd_sc_hd__buf_4 _0781_ (.A(_0088_),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_8 _0782_ (.A(_0094_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2i_1 _0783_ (.A0(\active_row[4][12] ),
    .A1(\active_row[6][12] ),
    .S(_0107_),
    .Y(_0143_));
 sky130_fd_sc_hd__nand3b_1 _0784_ (.A_N(_0121_),
    .B(\active_row[5][12] ),
    .C(_0142_),
    .Y(_0144_));
 sky130_fd_sc_hd__o21ai_0 _0785_ (.A1(_0142_),
    .A2(_0143_),
    .B1(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__mux2i_1 _0786_ (.A0(\active_row[3][12] ),
    .A1(\active_row[7][12] ),
    .S(_0141_),
    .Y(_0146_));
 sky130_fd_sc_hd__nor3_1 _0787_ (.A(_0105_),
    .B(_0101_),
    .C(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__nor2b_1 _0788_ (.A(_0092_),
    .B_N(\active_row[1][12] ),
    .Y(_0148_));
 sky130_fd_sc_hd__o221a_1 _0789_ (.A1(_0101_),
    .A2(\active_row[2][12] ),
    .B1(_0148_),
    .B2(_0105_),
    .C1(_0104_),
    .X(_0149_));
 sky130_fd_sc_hd__a211oi_1 _0790_ (.A1(_0141_),
    .A2(_0145_),
    .B1(_0147_),
    .C1(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _0791_ (.A(\active_row[0][12] ),
    .B(_0114_),
    .Y(_0151_));
 sky130_fd_sc_hd__or3_1 _0792_ (.A(net18),
    .B(_0150_),
    .C(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__o21ai_0 _0793_ (.A1(_0150_),
    .A2(_0151_),
    .B1(net18),
    .Y(_0153_));
 sky130_fd_sc_hd__nand4_1 _0794_ (.A(_0139_),
    .B(_0140_),
    .C(_0152_),
    .D(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__mux2i_1 _0795_ (.A0(\active_row[6][11] ),
    .A1(\active_row[7][11] ),
    .S(_0142_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_1 _0796_ (.A(_0096_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21ai_0 _0797_ (.A1(_0101_),
    .A2(\active_row[2][11] ),
    .B1(_0134_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_1 _0798_ (.A(\active_row[4][11] ),
    .B(_0135_),
    .Y(_0158_));
 sky130_fd_sc_hd__mux2i_1 _0799_ (.A0(\active_row[1][11] ),
    .A1(\active_row[5][11] ),
    .S(_0088_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _0800_ (.A(_0107_),
    .B(\active_row[3][11] ),
    .Y(_0160_));
 sky130_fd_sc_hd__o32a_1 _0801_ (.A1(_0105_),
    .A2(_0092_),
    .A3(_0159_),
    .B1(_0160_),
    .B2(_0111_),
    .X(_0161_));
 sky130_fd_sc_hd__and4b_1 _0802_ (.A_N(_0156_),
    .B(_0157_),
    .C(_0158_),
    .D(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_1 _0803_ (.A(\active_row[0][8] ),
    .Y(_0163_));
 sky130_fd_sc_hd__nor3_1 _0804_ (.A(_0087_),
    .B(_0093_),
    .C(_0090_),
    .Y(_0164_));
 sky130_fd_sc_hd__a21oi_1 _0805_ (.A1(_0163_),
    .A2(_0164_),
    .B1(net14),
    .Y(_0165_));
 sky130_fd_sc_hd__mux2i_1 _0806_ (.A0(\active_row[5][8] ),
    .A1(\active_row[7][8] ),
    .S(_0089_),
    .Y(_0166_));
 sky130_fd_sc_hd__a21oi_1 _0807_ (.A1(_0089_),
    .A2(\active_row[6][8] ),
    .B1(net3),
    .Y(_0167_));
 sky130_fd_sc_hd__a211oi_1 _0808_ (.A1(_0093_),
    .A2(_0166_),
    .B1(_0167_),
    .C1(_0103_),
    .Y(_0168_));
 sky130_fd_sc_hd__mux2i_1 _0809_ (.A0(\active_row[1][8] ),
    .A1(\active_row[3][8] ),
    .S(_0089_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _0810_ (.A(_0111_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__o21a_1 _0811_ (.A1(_0100_),
    .A2(\active_row[2][8] ),
    .B1(_0134_),
    .X(_0171_));
 sky130_fd_sc_hd__a2111oi_2 _0812_ (.A1(\active_row[4][8] ),
    .A2(_0135_),
    .B1(_0168_),
    .C1(_0170_),
    .D1(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(_0165_),
    .A1(net14),
    .S(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2i_1 _0814_ (.A0(\active_row[1][10] ),
    .A1(\active_row[3][10] ),
    .S(_0090_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand3b_1 _0815_ (.A_N(_0091_),
    .B(\active_row[5][10] ),
    .C(_0087_),
    .Y(_0175_));
 sky130_fd_sc_hd__o21ai_0 _0816_ (.A1(_0088_),
    .A2(_0174_),
    .B1(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand2b_1 _0817_ (.A_N(\active_row[2][10] ),
    .B(_0090_),
    .Y(_0177_));
 sky130_fd_sc_hd__mux2_1 _0818_ (.A0(\active_row[6][10] ),
    .A1(\active_row[7][10] ),
    .S(_0093_),
    .X(_0178_));
 sky130_fd_sc_hd__a222oi_1 _0819_ (.A1(\active_row[4][10] ),
    .A2(_0135_),
    .B1(_0177_),
    .B2(_0134_),
    .C1(_0178_),
    .C2(_0131_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21boi_2 _0820_ (.A1(_0097_),
    .A2(_0176_),
    .B1_N(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_1 _0821_ (.A(net16),
    .Y(_0181_));
 sky130_fd_sc_hd__o21ai_0 _0822_ (.A1(\active_row[0][10] ),
    .A2(_0113_),
    .B1(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(_0180_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(\active_row[1][6] ),
    .A1(\active_row[3][6] ),
    .S(_0092_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2b_1 _0825_ (.A_N(_0097_),
    .B(_0092_),
    .Y(_0185_));
 sky130_fd_sc_hd__o22ai_1 _0826_ (.A1(_0105_),
    .A2(_0184_),
    .B1(_0185_),
    .B2(\active_row[2][6] ),
    .Y(_0186_));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(\active_row[0][6] ),
    .B(_0114_),
    .Y(_0187_));
 sky130_fd_sc_hd__mux4_1 _0828_ (.A0(\active_row[4][6] ),
    .A1(\active_row[5][6] ),
    .A2(\active_row[6][6] ),
    .A3(\active_row[7][6] ),
    .S0(_0097_),
    .S1(_0121_),
    .X(_0188_));
 sky130_fd_sc_hd__nand3b_1 _0829_ (.A_N(net12),
    .B(_0188_),
    .C(_0141_),
    .Y(_0189_));
 sky130_fd_sc_hd__o41ai_1 _0830_ (.A1(_0141_),
    .A2(net12),
    .A3(_0186_),
    .A4(_0187_),
    .B1(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__o211ai_1 _0831_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0104_),
    .C1(net12),
    .Y(_0191_));
 sky130_fd_sc_hd__nand3b_1 _0832_ (.A_N(_0188_),
    .B(net12),
    .C(_0141_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand3b_1 _0833_ (.A_N(_0190_),
    .B(_0191_),
    .C(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__a2111o_1 _0834_ (.A1(net17),
    .A2(_0162_),
    .B1(_0173_),
    .C1(_0183_),
    .D1(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__o21ai_0 _0835_ (.A1(\active_row[0][7] ),
    .A2(_0114_),
    .B1(net13),
    .Y(_0195_));
 sky130_fd_sc_hd__mux2i_1 _0836_ (.A0(\active_row[1][7] ),
    .A1(\active_row[3][7] ),
    .S(_0107_),
    .Y(_0196_));
 sky130_fd_sc_hd__a2bb2oi_1 _0837_ (.A1_N(\active_row[2][7] ),
    .A2_N(_0185_),
    .B1(_0196_),
    .B2(_0142_),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(net13),
    .A1(_0195_),
    .S(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__mux4_1 _0839_ (.A0(\active_row[4][7] ),
    .A1(\active_row[5][7] ),
    .A2(\active_row[6][7] ),
    .A3(\active_row[7][7] ),
    .S0(_0097_),
    .S1(_0121_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0840_ (.A(net13),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor3_1 _0841_ (.A(\active_row[0][7] ),
    .B(net13),
    .C(_0114_),
    .Y(_0201_));
 sky130_fd_sc_hd__a21oi_1 _0842_ (.A1(_0141_),
    .A2(_0200_),
    .B1(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__o21ai_1 _0843_ (.A1(_0141_),
    .A2(_0198_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_1 _0844_ (.A(\active_row[5][4] ),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _0845_ (.A(_0121_),
    .B(\active_row[3][4] ),
    .Y(_0205_));
 sky130_fd_sc_hd__o32ai_4 _0846_ (.A1(_0107_),
    .A2(_0204_),
    .A3(_0109_),
    .B1(_0205_),
    .B2(_0111_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2b_1 _0847_ (.A(_0093_),
    .B_N(_0087_),
    .Y(_0207_));
 sky130_fd_sc_hd__nor4bb_1 _0848_ (.A(_0087_),
    .B(_0091_),
    .C_N(\active_row[1][4] ),
    .D_N(_0094_),
    .Y(_0208_));
 sky130_fd_sc_hd__a31o_1 _0849_ (.A1(_0101_),
    .A2(\active_row[4][4] ),
    .A3(_0207_),
    .B1(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2b_1 _0850_ (.A(\active_row[2][4] ),
    .B_N(_0092_),
    .Y(_0210_));
 sky130_fd_sc_hd__mux2i_1 _0851_ (.A0(\active_row[6][4] ),
    .A1(\active_row[7][4] ),
    .S(_0142_),
    .Y(_0211_));
 sky130_fd_sc_hd__o32ai_2 _0852_ (.A1(_0141_),
    .A2(_0142_),
    .A3(_0210_),
    .B1(_0211_),
    .B2(_0096_),
    .Y(_0212_));
 sky130_fd_sc_hd__o32ai_4 _0853_ (.A1(_0206_),
    .A2(_0209_),
    .A3(_0212_),
    .B1(_0114_),
    .B2(\active_row[0][4] ),
    .Y(_0213_));
 sky130_fd_sc_hd__xor2_1 _0854_ (.A(net9),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _0855_ (.A(_0203_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor4_2 _0856_ (.A(_0127_),
    .B(_0154_),
    .C(_0194_),
    .D(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_1 _0857_ (.A(\active_row[0][11] ),
    .Y(_0217_));
 sky130_fd_sc_hd__a211oi_1 _0858_ (.A1(_0217_),
    .A2(_0164_),
    .B1(_0162_),
    .C1(net17),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_1 _0859_ (.A(net6),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_1 _0860_ (.A(\active_row[5][1] ),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _0861_ (.A(_0121_),
    .B(\active_row[3][1] ),
    .Y(_0221_));
 sky130_fd_sc_hd__o32ai_2 _0862_ (.A1(_0121_),
    .A2(_0220_),
    .A3(_0109_),
    .B1(_0221_),
    .B2(_0111_),
    .Y(_0222_));
 sky130_fd_sc_hd__nor4bb_1 _0863_ (.A(_0088_),
    .B(_0092_),
    .C_N(\active_row[1][1] ),
    .D_N(_0097_),
    .Y(_0223_));
 sky130_fd_sc_hd__a31o_1 _0864_ (.A1(_0101_),
    .A2(\active_row[4][1] ),
    .A3(_0207_),
    .B1(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__nor2b_1 _0865_ (.A(\active_row[2][1] ),
    .B_N(_0107_),
    .Y(_0225_));
 sky130_fd_sc_hd__mux2i_2 _0866_ (.A0(\active_row[6][1] ),
    .A1(\active_row[7][1] ),
    .S(_0142_),
    .Y(_0226_));
 sky130_fd_sc_hd__o32ai_4 _0867_ (.A1(_0141_),
    .A2(_0142_),
    .A3(_0225_),
    .B1(_0226_),
    .B2(_0096_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor4_1 _0868_ (.A(_0219_),
    .B(_0222_),
    .C(_0224_),
    .D(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor3_1 _0869_ (.A(_0222_),
    .B(_0224_),
    .C(_0227_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_0 _0870_ (.A1(\active_row[0][1] ),
    .A2(_0114_),
    .B1(_0219_),
    .Y(_0230_));
 sky130_fd_sc_hd__o2bb2ai_1 _0871_ (.A1_N(net16),
    .A2_N(_0180_),
    .B1(_0229_),
    .B2(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__or3_1 _0872_ (.A(_0218_),
    .B(_0228_),
    .C(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__nand2_1 _0873_ (.A(_0107_),
    .B(\active_row[3][0] ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand3b_1 _0874_ (.A_N(_0092_),
    .B(\active_row[5][0] ),
    .C(_0088_),
    .Y(_0234_));
 sky130_fd_sc_hd__o21ai_0 _0875_ (.A1(_0088_),
    .A2(_0233_),
    .B1(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2b_1 _0876_ (.A_N(\active_row[1][0] ),
    .B(_0094_),
    .Y(_0236_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(_0105_),
    .A2(\active_row[4][0] ),
    .B1(_0236_),
    .B2(_0104_),
    .X(_0237_));
 sky130_fd_sc_hd__a22oi_1 _0878_ (.A1(_0142_),
    .A2(_0235_),
    .B1(_0237_),
    .B2(_0101_),
    .Y(_0238_));
 sky130_fd_sc_hd__mux2i_1 _0879_ (.A0(\active_row[6][0] ),
    .A1(\active_row[7][0] ),
    .S(_0097_),
    .Y(_0239_));
 sky130_fd_sc_hd__o2bb2ai_1 _0880_ (.A1_N(\active_row[2][0] ),
    .A2_N(_0134_),
    .B1(_0239_),
    .B2(_0104_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(_0121_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__o2bb2ai_1 _0882_ (.A1_N(_0238_),
    .A2_N(_0241_),
    .B1(_0114_),
    .B2(\active_row[0][0] ),
    .Y(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0883_ (.A(net5),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_1 _0884_ (.A(\active_row[0][13] ),
    .Y(_0244_));
 sky130_fd_sc_hd__a222oi_1 _0885_ (.A1(_0163_),
    .A2(net14),
    .B1(_0217_),
    .B2(net17),
    .C1(_0244_),
    .C2(net19),
    .Y(_0245_));
 sky130_fd_sc_hd__o221ai_1 _0886_ (.A1(\active_row[0][1] ),
    .A2(_0219_),
    .B1(\active_row[0][10] ),
    .B2(_0181_),
    .C1(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__mux4_1 _0887_ (.A0(\bank_active[0] ),
    .A1(\bank_active[1] ),
    .A2(\bank_active[2] ),
    .A3(\bank_active[3] ),
    .S0(_0094_),
    .S1(_0107_),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(_0141_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__mux4_1 _0889_ (.A0(\bank_active[4] ),
    .A1(\bank_active[5] ),
    .A2(\bank_active[6] ),
    .A3(\bank_active[7] ),
    .S0(_0094_),
    .S1(_0107_),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _0890_ (.A(_0104_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__a211o_1 _0891_ (.A1(net7),
    .A2(_0138_),
    .B1(_0248_),
    .C1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__a21oi_1 _0892_ (.A1(_0164_),
    .A2(_0246_),
    .B1(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__mux2_1 _0893_ (.A0(\active_row[1][13] ),
    .A1(\active_row[3][13] ),
    .S(_0090_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2i_2 _0894_ (.A0(\active_row[4][13] ),
    .A1(\active_row[6][13] ),
    .S(_0091_),
    .Y(_0254_));
 sky130_fd_sc_hd__a2bb2oi_1 _0895_ (.A1_N(_0111_),
    .A2_N(_0253_),
    .B1(_0254_),
    .B2(_0207_),
    .Y(_0255_));
 sky130_fd_sc_hd__mux2i_1 _0896_ (.A0(\active_row[5][13] ),
    .A1(\active_row[7][13] ),
    .S(_0091_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor4b_1 _0897_ (.A(_0087_),
    .B(_0094_),
    .C(\active_row[2][13] ),
    .D_N(_0091_),
    .Y(_0257_));
 sky130_fd_sc_hd__a31oi_1 _0898_ (.A1(_0088_),
    .A2(_0097_),
    .A3(_0256_),
    .B1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_1 _0899_ (.A(net19),
    .Y(_0259_));
 sky130_fd_sc_hd__o2111ai_1 _0900_ (.A1(\active_row[0][13] ),
    .A2(_0113_),
    .B1(_0255_),
    .C1(_0258_),
    .D1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _0901_ (.A(_0255_),
    .B(_0258_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _0902_ (.A(net19),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand3_1 _0903_ (.A(_0252_),
    .B(_0260_),
    .C(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nor3_2 _0904_ (.A(_0232_),
    .B(_0243_),
    .C(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2b_1 _0905_ (.A(_0090_),
    .B_N(\active_row[4][5] ),
    .Y(_0265_));
 sky130_fd_sc_hd__a211oi_1 _0906_ (.A1(_0091_),
    .A2(\active_row[6][5] ),
    .B1(_0265_),
    .C1(_0094_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0907_ (.A1(_0100_),
    .A2(\active_row[5][5] ),
    .B1(_0105_),
    .Y(_0267_));
 sky130_fd_sc_hd__mux2i_1 _0908_ (.A0(\active_row[2][5] ),
    .A1(\active_row[3][5] ),
    .S(_0093_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21boi_0 _0909_ (.A1(_0094_),
    .A2(\active_row[7][5] ),
    .B1_N(_0087_),
    .Y(_0269_));
 sky130_fd_sc_hd__a211o_1 _0910_ (.A1(_0103_),
    .A2(_0268_),
    .B1(_0269_),
    .C1(_0101_),
    .X(_0270_));
 sky130_fd_sc_hd__o211ai_1 _0911_ (.A1(_0105_),
    .A2(\active_row[1][5] ),
    .B1(_0101_),
    .C1(_0104_),
    .Y(_0271_));
 sky130_fd_sc_hd__o311a_1 _0912_ (.A1(_0104_),
    .A2(_0266_),
    .A3(_0267_),
    .B1(_0270_),
    .C1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _0913_ (.A(\active_row[0][5] ),
    .B(_0114_),
    .Y(_0273_));
 sky130_fd_sc_hd__or3_1 _0914_ (.A(net10),
    .B(_0272_),
    .C(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_0 _0915_ (.A1(_0272_),
    .A2(_0273_),
    .B1(net10),
    .Y(_0275_));
 sky130_fd_sc_hd__and2_1 _0916_ (.A(_0274_),
    .B(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _0917_ (.A(net32),
    .B(_0053_),
    .C(_0057_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _0918_ (.A(net33),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_1 _0919_ (.A(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand4_4 _0920_ (.A(_0216_),
    .B(_0264_),
    .C(_0276_),
    .D(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _0921_ (.A(_0664_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _0922_ (.A(\refresh_counter[15] ),
    .B(\refresh_counter[14] ),
    .C(\refresh_counter[13] ),
    .D(\refresh_counter[12] ),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_1 _0923_ (.A(\refresh_counter[6] ),
    .B(\refresh_counter[5] ),
    .Y(_0283_));
 sky130_fd_sc_hd__o2111ai_1 _0924_ (.A1(_0645_),
    .A2(_0643_),
    .B1(\refresh_counter[4] ),
    .C1(\refresh_counter[3] ),
    .D1(\refresh_counter[2] ),
    .Y(_0284_));
 sky130_fd_sc_hd__nand4_1 _0925_ (.A(\refresh_counter[10] ),
    .B(\refresh_counter[9] ),
    .C(\refresh_counter[8] ),
    .D(\refresh_counter[7] ),
    .Y(_0285_));
 sky130_fd_sc_hd__a21oi_1 _0926_ (.A1(_0283_),
    .A2(_0284_),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__or3_1 _0927_ (.A(\refresh_counter[11] ),
    .B(_0282_),
    .C(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_4 _0928_ (.A(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _0929_ (.A(_0288_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_2 _0930_ (.A(_0281_),
    .B(_0639_),
    .Y(_0289_));
 sky130_fd_sc_hd__clkbuf_4 _0931_ (.A(_0083_),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_4 _0932_ (.A(_0070_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _0933_ (.A(_0291_),
    .B(net33),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_1 _0934_ (.A(\burst_counter[2] ),
    .B(\burst_counter[3] ),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_2 _0935_ (.A(_0635_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand4b_1 _0936_ (.A_N(net133),
    .B(_0086_),
    .C(_0294_),
    .D(_0084_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_0 _0937_ (.A1(_0290_),
    .A2(_0292_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__a2bb2oi_1 _0938_ (.A1_N(_0280_),
    .A2_N(_0289_),
    .B1(_0296_),
    .B2(_0067_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _0939_ (.A(_0062_),
    .B(_0297_),
    .Y(_0670_));
 sky130_fd_sc_hd__clkinv_2 _0940_ (.A(_0664_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _0941_ (.A(_0280_),
    .B(_0288_),
    .Y(_0299_));
 sky130_fd_sc_hd__clkinvlp_4 _0942_ (.A(_0070_),
    .Y(_0300_));
 sky130_fd_sc_hd__a21oi_1 _0943_ (.A1(net33),
    .A2(_0067_),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nor2_2 _0944_ (.A(_0050_),
    .B(_0070_),
    .Y(_0302_));
 sky130_fd_sc_hd__nor2_1 _0945_ (.A(_0664_),
    .B(_0083_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_4 _0946_ (.A(_0302_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_1 _0947_ (.A(_0065_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21ai_4 _0948_ (.A1(_0305_),
    .A2(_0294_),
    .B1(_0083_),
    .Y(_0306_));
 sky130_fd_sc_hd__buf_2 _0949_ (.A(_0305_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_2 _0950_ (.A(_0072_),
    .B(\init_state[1] ),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _0951_ (.A(\init_state[6] ),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__o21ai_2 _0952_ (.A1(_0307_),
    .A2(_0309_),
    .B1(_0050_),
    .Y(_0310_));
 sky130_fd_sc_hd__nand3_1 _0953_ (.A(_0304_),
    .B(_0306_),
    .C(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_1 _0954_ (.A(_0301_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__o21ai_1 _0955_ (.A1(_0298_),
    .A2(_0299_),
    .B1(_0312_),
    .Y(_0583_));
 sky130_fd_sc_hd__o21ai_4 _0956_ (.A1(_0063_),
    .A2(_0064_),
    .B1(_0070_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21boi_0 _0957_ (.A1(_0300_),
    .A2(_0298_),
    .B1_N(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__o21ai_0 _0958_ (.A1(_0062_),
    .A2(_0314_),
    .B1(_0310_),
    .Y(_0315_));
 sky130_fd_sc_hd__nor2_1 _0959_ (.A(_0085_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand3_2 _0960_ (.A(net32),
    .B(_0053_),
    .C(_0057_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand3_4 _0961_ (.A(_0216_),
    .B(_0264_),
    .C(_0276_),
    .Y(_0318_));
 sky130_fd_sc_hd__buf_4 _0962_ (.A(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_4 _0963_ (.A(_0298_),
    .B(_0288_),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_0 _0964_ (.A1(_0317_),
    .A2(_0319_),
    .B1(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _0965_ (.A(_0316_),
    .B(_0321_),
    .Y(_0584_));
 sky130_fd_sc_hd__a21oi_1 _0966_ (.A1(_0277_),
    .A2(_0318_),
    .B1(_0289_),
    .Y(_0322_));
 sky130_fd_sc_hd__or3_1 _0967_ (.A(_0291_),
    .B(_0311_),
    .C(_0322_),
    .X(_0585_));
 sky130_fd_sc_hd__nor2_2 _0968_ (.A(_0050_),
    .B(_0281_),
    .Y(_0323_));
 sky130_fd_sc_hd__a21boi_4 _0969_ (.A1(\init_state[7] ),
    .A2(_0066_),
    .B1_N(_0050_),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_1 _0970_ (.A(_0323_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__clkbuf_4 _0971_ (.A(_0281_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0972_ (.A(_0326_),
    .B(_0641_),
    .Y(_0327_));
 sky130_fd_sc_hd__o21ai_0 _0973_ (.A1(_0642_),
    .A2(_0325_),
    .B1(_0327_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor3_4 _0974_ (.A(_0320_),
    .B(_0323_),
    .C(_0324_),
    .Y(_0328_));
 sky130_fd_sc_hd__buf_2 _0975_ (.A(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _0976_ (.A(\refresh_counter[1] ),
    .B(_0639_),
    .Y(_0330_));
 sky130_fd_sc_hd__a211oi_1 _0977_ (.A1(_0644_),
    .A2(_0639_),
    .B1(_0329_),
    .C1(_0330_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _0978_ (.A(_0645_),
    .B(_0639_),
    .Y(_0331_));
 sky130_fd_sc_hd__xor2_1 _0979_ (.A(\refresh_counter[2] ),
    .B(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(_0329_),
    .B(_0332_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand4_1 _0981_ (.A(\refresh_counter[2] ),
    .B(\refresh_counter[1] ),
    .C(\refresh_counter[0] ),
    .D(_0639_),
    .Y(_0333_));
 sky130_fd_sc_hd__xor2_1 _0982_ (.A(\refresh_counter[3] ),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_1 _0983_ (.A(_0329_),
    .B(_0334_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand4_1 _0984_ (.A(\refresh_counter[3] ),
    .B(\refresh_counter[2] ),
    .C(_0645_),
    .D(_0639_),
    .Y(_0335_));
 sky130_fd_sc_hd__xor2_1 _0985_ (.A(\refresh_counter[4] ),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(_0329_),
    .B(_0336_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(\refresh_counter[4] ),
    .B(\refresh_counter[3] ),
    .Y(_0337_));
 sky130_fd_sc_hd__nor2_1 _0988_ (.A(_0337_),
    .B(_0333_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_1 _0989_ (.A(\refresh_counter[5] ),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nor2_1 _0990_ (.A(_0329_),
    .B(_0339_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand3_1 _0991_ (.A(\refresh_counter[4] ),
    .B(\refresh_counter[3] ),
    .C(\refresh_counter[2] ),
    .Y(_0340_));
 sky130_fd_sc_hd__nor2_1 _0992_ (.A(_0340_),
    .B(_0331_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(\refresh_counter[5] ),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__xor2_1 _0994_ (.A(\refresh_counter[6] ),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_1 _0995_ (.A(_0329_),
    .B(_0343_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3_1 _0996_ (.A(\refresh_counter[6] ),
    .B(\refresh_counter[5] ),
    .C(_0338_),
    .Y(_0344_));
 sky130_fd_sc_hd__xor2_1 _0997_ (.A(\refresh_counter[7] ),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__nor2_1 _0998_ (.A(_0329_),
    .B(_0345_),
    .Y(_0599_));
 sky130_fd_sc_hd__and3_1 _0999_ (.A(\refresh_counter[7] ),
    .B(\refresh_counter[6] ),
    .C(\refresh_counter[5] ),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _1000_ (.A(_0341_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__xor2_1 _1001_ (.A(\refresh_counter[8] ),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(_0329_),
    .B(_0348_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand3_1 _1003_ (.A(\refresh_counter[8] ),
    .B(_0338_),
    .C(_0346_),
    .Y(_0349_));
 sky130_fd_sc_hd__xor2_1 _1004_ (.A(\refresh_counter[9] ),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(_0329_),
    .B(_0350_),
    .Y(_0601_));
 sky130_fd_sc_hd__a41oi_1 _1006_ (.A1(\refresh_counter[9] ),
    .A2(\refresh_counter[8] ),
    .A3(_0341_),
    .A4(_0346_),
    .B1(\refresh_counter[10] ),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_1 _1007_ (.A(_0329_),
    .B(_0351_),
    .Y(_0587_));
 sky130_fd_sc_hd__nor2b_1 _1008_ (.A(_0328_),
    .B_N(\refresh_counter[11] ),
    .Y(_0588_));
 sky130_fd_sc_hd__nor2b_1 _1009_ (.A(_0328_),
    .B_N(\refresh_counter[12] ),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2b_1 _1010_ (.A(_0328_),
    .B_N(\refresh_counter[13] ),
    .Y(_0590_));
 sky130_fd_sc_hd__nor2b_1 _1011_ (.A(_0328_),
    .B_N(\refresh_counter[14] ),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2b_1 _1012_ (.A(_0328_),
    .B_N(\refresh_counter[15] ),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_1 _1013_ (.A(\timer[0] ),
    .Y(_0647_));
 sky130_fd_sc_hd__or2_0 _1014_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(net133),
    .B(_0086_),
    .Y(_0353_));
 sky130_fd_sc_hd__nor3_2 _1016_ (.A(_0352_),
    .B(_0064_),
    .C(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nor3_1 _1017_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[1] ),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_1 _1018_ (.A(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__o21ai_0 _1019_ (.A1(_0656_),
    .A2(_0356_),
    .B1(_0354_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2b_1 _1020_ (.A_N(net133),
    .B(net101),
    .Y(_0358_));
 sky130_fd_sc_hd__nand3_1 _1021_ (.A(net133),
    .B(net198),
    .C(net35),
    .Y(_0359_));
 sky130_fd_sc_hd__a21boi_1 _1022_ (.A1(_0358_),
    .A2(_0359_),
    .B1_N(_0086_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _1023_ (.A(_0294_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__o21ai_0 _1024_ (.A1(_0650_),
    .A2(_0360_),
    .B1(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a32oi_1 _1025_ (.A1(_0647_),
    .A2(_0354_),
    .A3(_0356_),
    .B1(_0357_),
    .B2(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_1 _1026_ (.A(_0650_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand3_1 _1027_ (.A(_0364_),
    .B(_0066_),
    .C(_0294_),
    .Y(_0365_));
 sky130_fd_sc_hd__o21ai_0 _1028_ (.A1(_0066_),
    .A2(_0363_),
    .B1(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nor3_2 _1029_ (.A(\init_state[2] ),
    .B(\init_state[6] ),
    .C(_0308_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor3_1 _1030_ (.A(\init_state[4] ),
    .B(\init_state[3] ),
    .C(\init_state[0] ),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(_0367_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(_0649_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__o21ai_0 _1033_ (.A1(_0650_),
    .A2(_0369_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__o21ai_0 _1034_ (.A1(_0300_),
    .A2(_0651_),
    .B1(_0304_),
    .Y(_0372_));
 sky130_fd_sc_hd__a221o_1 _1035_ (.A1(_0083_),
    .A2(_0366_),
    .B1(_0371_),
    .B2(_0061_),
    .C1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__o21a_1 _1036_ (.A1(_0277_),
    .A2(_0373_),
    .B1(_0304_),
    .X(_0374_));
 sky130_fd_sc_hd__o22a_1 _1037_ (.A1(_0322_),
    .A2(_0373_),
    .B1(_0374_),
    .B2(_0364_),
    .X(_0602_));
 sky130_fd_sc_hd__inv_1 _1038_ (.A(\timer[1] ),
    .Y(_0653_));
 sky130_fd_sc_hd__clkbuf_4 _1039_ (.A(_0307_),
    .X(_0648_));
 sky130_fd_sc_hd__a211oi_1 _1040_ (.A1(net32),
    .A2(_0304_),
    .B1(_0307_),
    .C1(\timer[1] ),
    .Y(_0375_));
 sky130_fd_sc_hd__a21oi_1 _1041_ (.A1(_0655_),
    .A2(_0648_),
    .B1(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__and2_2 _1042_ (.A(_0635_),
    .B(_0293_),
    .X(_0377_));
 sky130_fd_sc_hd__nor4_1 _1043_ (.A(_0352_),
    .B(_0054_),
    .C(_0055_),
    .D(_0056_),
    .Y(_0378_));
 sky130_fd_sc_hd__a41oi_1 _1044_ (.A1(net133),
    .A2(_0656_),
    .A3(_0086_),
    .A4(_0378_),
    .B1(_0360_),
    .Y(_0379_));
 sky130_fd_sc_hd__a21oi_2 _1045_ (.A1(_0354_),
    .A2(_0356_),
    .B1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_0 _1046_ (.A1(_0655_),
    .A2(_0380_),
    .B1(_0307_),
    .Y(_0381_));
 sky130_fd_sc_hd__o311ai_0 _1047_ (.A1(\timer[1] ),
    .A2(_0307_),
    .A3(_0377_),
    .B1(_0381_),
    .C1(_0083_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(\timer[1] ),
    .B(_0368_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _1049_ (.A(_0066_),
    .B(_0367_),
    .C(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21o_1 _1050_ (.A1(net33),
    .A2(_0066_),
    .B1(_0300_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _1051_ (.A(_0385_),
    .B(_0304_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _1052_ (.A1(_0061_),
    .A2(_0384_),
    .B1(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor3_1 _1053_ (.A(\timer[1] ),
    .B(_0307_),
    .C(_0304_),
    .Y(_0388_));
 sky130_fd_sc_hd__a221oi_1 _1054_ (.A1(_0655_),
    .A2(_0307_),
    .B1(_0382_),
    .B2(_0387_),
    .C1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__a31o_1 _1055_ (.A1(_0280_),
    .A2(_0320_),
    .A3(_0376_),
    .B1(_0389_),
    .X(_0609_));
 sky130_fd_sc_hd__xor2_1 _1056_ (.A(\timer[2] ),
    .B(_0654_),
    .X(_0390_));
 sky130_fd_sc_hd__a21oi_1 _1057_ (.A1(_0307_),
    .A2(_0390_),
    .B1(_0288_),
    .Y(_0391_));
 sky130_fd_sc_hd__o31ai_1 _1058_ (.A1(net33),
    .A2(_0317_),
    .A3(_0318_),
    .B1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_0 _1059_ (.A1(_0307_),
    .A2(_0301_),
    .B1(_0390_),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2b_1 _1060_ (.A(_0380_),
    .B_N(_0083_),
    .Y(_0394_));
 sky130_fd_sc_hd__nor3_1 _1061_ (.A(_0061_),
    .B(_0386_),
    .C(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _1062_ (.A1(_0075_),
    .A2(_0393_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a21o_1 _1063_ (.A1(_0326_),
    .A2(_0392_),
    .B1(_0396_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(\init_state[4] ),
    .B(\init_state[3] ),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _1065_ (.A(_0367_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__a221oi_1 _1066_ (.A1(_0290_),
    .A2(_0377_),
    .B1(_0398_),
    .B2(_0062_),
    .C1(_0648_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand4_1 _1067_ (.A(net32),
    .B(_0280_),
    .C(_0320_),
    .D(_0304_),
    .Y(_0400_));
 sky130_fd_sc_hd__nor3_1 _1068_ (.A(\timer[2] ),
    .B(\timer[1] ),
    .C(\timer[0] ),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_1 _1069_ (.A(\timer[3] ),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__nor2_1 _1070_ (.A(_0289_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nor2_1 _1071_ (.A(_0395_),
    .B(_0402_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor3_1 _1072_ (.A(_0067_),
    .B(_0403_),
    .C(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__a31oi_1 _1073_ (.A1(_0385_),
    .A2(_0399_),
    .A3(_0400_),
    .B1(_0405_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand2_1 _1074_ (.A(_0654_),
    .B(_0052_),
    .Y(_0406_));
 sky130_fd_sc_hd__xor2_1 _1075_ (.A(\timer[4] ),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__nor2_1 _1076_ (.A(_0067_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _1077_ (.A(_0288_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o221ai_2 _1078_ (.A1(_0281_),
    .A2(_0084_),
    .B1(_0306_),
    .B2(_0380_),
    .C1(_0302_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21oi_1 _1079_ (.A1(_0408_),
    .A2(_0410_),
    .B1(_0326_),
    .Y(_0411_));
 sky130_fd_sc_hd__nor2_1 _1080_ (.A(_0409_),
    .B(_0411_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand3_1 _1081_ (.A(_0653_),
    .B(_0647_),
    .C(_0052_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_1 _1082_ (.A(\timer[4] ),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__xor2_1 _1083_ (.A(\timer[5] ),
    .B(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _1084_ (.A(_0648_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nand3_1 _1085_ (.A(_0062_),
    .B(\init_state[0] ),
    .C(_0067_),
    .Y(_0416_));
 sky130_fd_sc_hd__nor2_1 _1086_ (.A(_0320_),
    .B(_0410_),
    .Y(_0417_));
 sky130_fd_sc_hd__a21oi_1 _1087_ (.A1(_0415_),
    .A2(_0416_),
    .B1(_0417_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_0 _1088_ (.A1(_0066_),
    .A2(_0367_),
    .B1(_0368_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _1089_ (.A(_0061_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(_0050_),
    .B(_0309_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2b_1 _1091_ (.A_N(\init_state[2] ),
    .B(_0368_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21ai_0 _1092_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0304_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21oi_1 _1093_ (.A1(_0307_),
    .A2(_0380_),
    .B1(_0306_),
    .Y(_0423_));
 sky130_fd_sc_hd__a211oi_2 _1094_ (.A1(_0317_),
    .A2(_0320_),
    .B1(_0422_),
    .C1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__a211oi_1 _1095_ (.A1(_0057_),
    .A2(_0419_),
    .B1(\timer[6] ),
    .C1(_0063_),
    .Y(_0425_));
 sky130_fd_sc_hd__a21oi_1 _1096_ (.A1(\timer[6] ),
    .A2(_0063_),
    .B1(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31oi_1 _1097_ (.A1(_0300_),
    .A2(_0419_),
    .A3(_0424_),
    .B1(_0426_),
    .Y(_0614_));
 sky130_fd_sc_hd__a21oi_1 _1098_ (.A1(_0062_),
    .A2(_0369_),
    .B1(_0291_),
    .Y(_0427_));
 sky130_fd_sc_hd__or3_1 _1099_ (.A(\timer[6] ),
    .B(_0352_),
    .C(_0412_),
    .X(_0428_));
 sky130_fd_sc_hd__xnor2_1 _1100_ (.A(\timer[7] ),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor3b_1 _1101_ (.A(_0397_),
    .B(_0648_),
    .C_N(_0062_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21oi_1 _1102_ (.A1(_0648_),
    .A2(_0429_),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_1 _1103_ (.A1(_0424_),
    .A2(_0427_),
    .B1(_0431_),
    .Y(_0615_));
 sky130_fd_sc_hd__o21a_1 _1104_ (.A1(_0067_),
    .A2(_0302_),
    .B1(_0424_),
    .X(_0432_));
 sky130_fd_sc_hd__nor4_1 _1105_ (.A(\timer[7] ),
    .B(\timer[6] ),
    .C(_0063_),
    .D(_0378_),
    .Y(_0433_));
 sky130_fd_sc_hd__xnor2_1 _1106_ (.A(\timer[8] ),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__nor2_1 _1107_ (.A(_0432_),
    .B(_0434_),
    .Y(_0616_));
 sky130_fd_sc_hd__nor3_1 _1108_ (.A(\timer[7] ),
    .B(\timer[8] ),
    .C(_0428_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _1109_ (.A(\timer[9] ),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _1110_ (.A(_0424_),
    .B(_0427_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_2 _1111_ (.A(_0648_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(_0436_),
    .B(_0438_),
    .Y(_0617_));
 sky130_fd_sc_hd__or3_1 _1113_ (.A(\timer[7] ),
    .B(\timer[9] ),
    .C(\timer[8] ),
    .X(_0439_));
 sky130_fd_sc_hd__nor3_1 _1114_ (.A(\timer[6] ),
    .B(_0063_),
    .C(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__xnor2_1 _1115_ (.A(\timer[10] ),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nor2_1 _1116_ (.A(_0438_),
    .B(_0441_),
    .Y(_0603_));
 sky130_fd_sc_hd__or3_1 _1117_ (.A(\timer[11] ),
    .B(_0054_),
    .C(_0428_),
    .X(_0442_));
 sky130_fd_sc_hd__o21ai_0 _1118_ (.A1(_0054_),
    .A2(_0428_),
    .B1(\timer[11] ),
    .Y(_0443_));
 sky130_fd_sc_hd__a21oi_1 _1119_ (.A1(_0442_),
    .A2(_0443_),
    .B1(_0438_),
    .Y(_0604_));
 sky130_fd_sc_hd__nor4b_1 _1120_ (.A(_0063_),
    .B(_0054_),
    .C(_0055_),
    .D_N(_0056_),
    .Y(_0444_));
 sky130_fd_sc_hd__xnor2_1 _1121_ (.A(\timer[12] ),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nor2_1 _1122_ (.A(_0432_),
    .B(_0445_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1123_ (.A(\timer[12] ),
    .B(_0442_),
    .Y(_0446_));
 sky130_fd_sc_hd__xnor2_1 _1124_ (.A(\timer[13] ),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _1125_ (.A(_0438_),
    .B(_0447_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _1127_ (.A(_0448_),
    .B(_0444_),
    .Y(_0449_));
 sky130_fd_sc_hd__xor2_1 _1128_ (.A(\timer[14] ),
    .B(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _1129_ (.A(_0432_),
    .B(_0450_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor4_1 _1130_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[14] ),
    .D(_0442_),
    .Y(_0451_));
 sky130_fd_sc_hd__xnor2_1 _1131_ (.A(\timer[15] ),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _1132_ (.A(_0438_),
    .B(_0452_),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_1 _1133_ (.A1(net35),
    .A2(_0294_),
    .B1(_0353_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _1134_ (.A(_0067_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand4_1 _1135_ (.A(_0656_),
    .B(_0648_),
    .C(_0354_),
    .D(_0355_),
    .Y(_0455_));
 sky130_fd_sc_hd__a21boi_0 _1136_ (.A1(_0454_),
    .A2(_0455_),
    .B1_N(_0085_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_1 _1137_ (.A(net118),
    .Y(_0618_));
 sky130_fd_sc_hd__inv_1 _1138_ (.A(\refresh_counter[0] ),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_1 _1139_ (.A(net199),
    .Y(_0658_));
 sky130_fd_sc_hd__inv_1 _1140_ (.A(net119),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_1 _1141_ (.A(\burst_counter[1] ),
    .Y(_0634_));
 sky130_fd_sc_hd__inv_1 _1142_ (.A(net200),
    .Y(_0659_));
 sky130_fd_sc_hd__mux2i_1 _1143_ (.A0(net2),
    .A1(net5),
    .S(_0318_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _1144_ (.A(_0061_),
    .B(_0308_),
    .Y(_0457_));
 sky130_fd_sc_hd__o21ai_1 _1145_ (.A1(_0317_),
    .A2(_0288_),
    .B1(_0664_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand4_4 _1146_ (.A(_0304_),
    .B(_0306_),
    .C(_0313_),
    .D(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2b_1 _1147_ (.A(_0459_),
    .B_N(_0310_),
    .Y(_0460_));
 sky130_fd_sc_hd__clkbuf_2 _1148_ (.A(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(net104),
    .A1(_0457_),
    .S(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0326_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__nor2_2 _1151_ (.A(_0061_),
    .B(_0459_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_1 _1152_ (.A1(_0308_),
    .A2(_0461_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a21o_1 _1153_ (.A1(_0291_),
    .A2(net2),
    .B1(_0290_),
    .X(_0466_));
 sky130_fd_sc_hd__o21ai_0 _1154_ (.A1(_0465_),
    .A2(_0466_),
    .B1(_0462_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_0 _1155_ (.A1(_0456_),
    .A2(_0463_),
    .B1(_0467_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand3_1 _1156_ (.A(_0281_),
    .B(_0319_),
    .C(_0464_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2b_1 _1157_ (.A_N(_0459_),
    .B(_0310_),
    .Y(_0469_));
 sky130_fd_sc_hd__buf_2 _1158_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__a22oi_1 _1159_ (.A1(net105),
    .A2(_0470_),
    .B1(_0464_),
    .B2(_0085_),
    .Y(_0471_));
 sky130_fd_sc_hd__o21ai_0 _1160_ (.A1(_0181_),
    .A2(_0468_),
    .B1(_0471_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand3_1 _1161_ (.A(_0326_),
    .B(net17),
    .C(_0319_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _1162_ (.A(\init_state[1] ),
    .B(_0066_),
    .Y(_0473_));
 sky130_fd_sc_hd__a21oi_2 _1163_ (.A1(_0061_),
    .A2(_0473_),
    .B1(_0459_),
    .Y(_0474_));
 sky130_fd_sc_hd__a21oi_1 _1164_ (.A1(_0061_),
    .A2(_0072_),
    .B1(_0083_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand4b_1 _1165_ (.A_N(_0072_),
    .B(\init_state[1] ),
    .C(_0461_),
    .D(_0062_),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_0 _1166_ (.A1(net106),
    .A2(_0461_),
    .B1(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a31oi_1 _1167_ (.A1(_0472_),
    .A2(_0474_),
    .A3(_0475_),
    .B1(_0477_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_1 _1168_ (.A(net18),
    .Y(_0478_));
 sky130_fd_sc_hd__a22oi_1 _1169_ (.A1(net107),
    .A2(_0470_),
    .B1(_0464_),
    .B2(_0085_),
    .Y(_0479_));
 sky130_fd_sc_hd__o21ai_0 _1170_ (.A1(_0478_),
    .A2(_0468_),
    .B1(_0479_),
    .Y(_0021_));
 sky130_fd_sc_hd__a22oi_1 _1171_ (.A1(net108),
    .A2(_0470_),
    .B1(_0464_),
    .B2(_0085_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_0 _1172_ (.A1(_0259_),
    .A2(_0468_),
    .B1(_0480_),
    .Y(_0022_));
 sky130_fd_sc_hd__mux2i_1 _1173_ (.A0(net11),
    .A1(net6),
    .S(_0318_),
    .Y(_0481_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(net109),
    .A1(_0457_),
    .S(_0461_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _1175_ (.A(_0326_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21o_1 _1176_ (.A1(_0291_),
    .A2(net11),
    .B1(_0290_),
    .X(_0484_));
 sky130_fd_sc_hd__o21ai_0 _1177_ (.A1(_0465_),
    .A2(_0484_),
    .B1(_0482_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21ai_0 _1178_ (.A1(_0481_),
    .A2(_0483_),
    .B1(_0485_),
    .Y(_0023_));
 sky130_fd_sc_hd__mux2i_1 _1179_ (.A0(net20),
    .A1(net7),
    .S(_0318_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0326_),
    .B(_0474_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_1 _1181_ (.A(_0050_),
    .B(_0083_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(_0291_),
    .B(net20),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _1183_ (.A(_0488_),
    .B(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__a22oi_1 _1184_ (.A1(net110),
    .A2(_0470_),
    .B1(_0474_),
    .B2(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_0 _1185_ (.A1(_0486_),
    .A2(_0487_),
    .B1(_0491_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(_0326_),
    .B(_0464_),
    .Y(_0492_));
 sky130_fd_sc_hd__mux2i_1 _1187_ (.A0(net21),
    .A1(net8),
    .S(_0319_),
    .Y(_0493_));
 sky130_fd_sc_hd__a21oi_1 _1188_ (.A1(_0291_),
    .A2(net21),
    .B1(_0290_),
    .Y(_0494_));
 sky130_fd_sc_hd__nor3_1 _1189_ (.A(_0062_),
    .B(_0459_),
    .C(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__a21oi_1 _1190_ (.A1(net111),
    .A2(_0470_),
    .B1(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__o21ai_0 _1191_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0496_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(_0072_),
    .B(_0066_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21oi_1 _1193_ (.A1(_0061_),
    .A2(_0497_),
    .B1(_0459_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_1 _1194_ (.A(_0281_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2i_1 _1195_ (.A0(net22),
    .A1(net9),
    .S(_0319_),
    .Y(_0500_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(_0070_),
    .A2(net22),
    .B1(_0059_),
    .B2(_0072_),
    .C1(_0084_),
    .X(_0501_));
 sky130_fd_sc_hd__a22oi_1 _1197_ (.A1(net112),
    .A2(_0470_),
    .B1(_0498_),
    .B2(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__o21ai_0 _1198_ (.A1(_0499_),
    .A2(_0500_),
    .B1(_0502_),
    .Y(_0026_));
 sky130_fd_sc_hd__mux2i_1 _1199_ (.A0(net23),
    .A1(net10),
    .S(_0318_),
    .Y(_0503_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(net113),
    .A1(_0457_),
    .S(_0461_),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _1201_ (.A(_0326_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a21o_1 _1202_ (.A1(_0291_),
    .A2(net23),
    .B1(_0290_),
    .X(_0506_));
 sky130_fd_sc_hd__o21ai_0 _1203_ (.A1(_0465_),
    .A2(_0506_),
    .B1(_0504_),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_0 _1204_ (.A1(_0503_),
    .A2(_0505_),
    .B1(_0507_),
    .Y(_0027_));
 sky130_fd_sc_hd__mux2i_1 _1205_ (.A0(net24),
    .A1(net12),
    .S(_0319_),
    .Y(_0508_));
 sky130_fd_sc_hd__a221o_1 _1206_ (.A1(_0070_),
    .A2(net24),
    .B1(_0058_),
    .B2(_0072_),
    .C1(_0084_),
    .X(_0509_));
 sky130_fd_sc_hd__a22oi_1 _1207_ (.A1(net114),
    .A2(_0470_),
    .B1(_0498_),
    .B2(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ai_0 _1208_ (.A1(_0499_),
    .A2(_0508_),
    .B1(_0510_),
    .Y(_0028_));
 sky130_fd_sc_hd__mux2i_1 _1209_ (.A0(net25),
    .A1(net13),
    .S(_0319_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21oi_1 _1210_ (.A1(_0291_),
    .A2(net25),
    .B1(_0290_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor3_1 _1211_ (.A(_0062_),
    .B(_0459_),
    .C(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__a21oi_1 _1212_ (.A1(net115),
    .A2(_0470_),
    .B1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o21ai_0 _1213_ (.A1(_0492_),
    .A2(_0511_),
    .B1(_0514_),
    .Y(_0029_));
 sky130_fd_sc_hd__mux2i_1 _1214_ (.A0(net26),
    .A1(net14),
    .S(_0319_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _1215_ (.A(_0291_),
    .B(net26),
    .Y(_0516_));
 sky130_fd_sc_hd__and3_1 _1216_ (.A(_0474_),
    .B(_0475_),
    .C(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__nand3_1 _1217_ (.A(_0474_),
    .B(_0475_),
    .C(_0516_),
    .Y(_0518_));
 sky130_fd_sc_hd__o221ai_1 _1218_ (.A1(net116),
    .A2(_0461_),
    .B1(_0518_),
    .B2(_0326_),
    .C1(_0476_),
    .Y(_0519_));
 sky130_fd_sc_hd__a21oi_1 _1219_ (.A1(_0515_),
    .A2(_0517_),
    .B1(_0519_),
    .Y(_0030_));
 sky130_fd_sc_hd__mux2i_1 _1220_ (.A0(net27),
    .A1(net15),
    .S(_0319_),
    .Y(_0520_));
 sky130_fd_sc_hd__a221o_1 _1221_ (.A1(_0070_),
    .A2(net27),
    .B1(_0058_),
    .B2(_0072_),
    .C1(_0084_),
    .X(_0521_));
 sky130_fd_sc_hd__a22oi_1 _1222_ (.A1(net117),
    .A2(_0470_),
    .B1(_0498_),
    .B2(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__o21ai_0 _1223_ (.A1(_0499_),
    .A2(_0520_),
    .B1(_0522_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand3_1 _1224_ (.A(_0084_),
    .B(_0377_),
    .C(_0323_),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_4 _1225_ (.A(_0648_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__and4b_1 _1226_ (.A_N(_0630_),
    .B(_0306_),
    .C(_0313_),
    .D(_0323_),
    .X(_0525_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(net120),
    .B(net119),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(net118),
    .B(_0621_),
    .Y(_0527_));
 sky130_fd_sc_hd__a31oi_1 _1229_ (.A1(_0525_),
    .A2(_0526_),
    .A3(_0527_),
    .B1(\bank_active[0] ),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(_0524_),
    .B(_0528_),
    .Y(_0032_));
 sky130_fd_sc_hd__and4_1 _1231_ (.A(_0630_),
    .B(_0306_),
    .C(_0313_),
    .D(_0323_),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _1232_ (.A1(_0624_),
    .A2(_0529_),
    .B1(\bank_active[1] ),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _1233_ (.A(_0524_),
    .B(_0530_),
    .Y(_0033_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(net118),
    .B(_0526_),
    .Y(_0531_));
 sky130_fd_sc_hd__a31oi_1 _1235_ (.A1(_0621_),
    .A2(_0529_),
    .A3(_0531_),
    .B1(\bank_active[2] ),
    .Y(_0532_));
 sky130_fd_sc_hd__nor2_1 _1236_ (.A(_0524_),
    .B(_0532_),
    .Y(_0034_));
 sky130_fd_sc_hd__a21oi_1 _1237_ (.A1(_0626_),
    .A2(_0529_),
    .B1(\bank_active[3] ),
    .Y(_0533_));
 sky130_fd_sc_hd__nor2_1 _1238_ (.A(_0524_),
    .B(_0533_),
    .Y(_0035_));
 sky130_fd_sc_hd__nor3_1 _1239_ (.A(net118),
    .B(_0621_),
    .C(_0526_),
    .Y(_0534_));
 sky130_fd_sc_hd__a21oi_1 _1240_ (.A1(_0529_),
    .A2(_0534_),
    .B1(\bank_active[4] ),
    .Y(_0535_));
 sky130_fd_sc_hd__nor2_1 _1241_ (.A(_0524_),
    .B(_0535_),
    .Y(_0036_));
 sky130_fd_sc_hd__a21oi_1 _1242_ (.A1(_0624_),
    .A2(_0525_),
    .B1(\bank_active[5] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(_0524_),
    .B(_0536_),
    .Y(_0037_));
 sky130_fd_sc_hd__a31oi_1 _1244_ (.A1(_0621_),
    .A2(_0525_),
    .A3(_0531_),
    .B1(\bank_active[6] ),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_1 _1245_ (.A(_0524_),
    .B(_0537_),
    .Y(_0038_));
 sky130_fd_sc_hd__a21oi_1 _1246_ (.A1(_0626_),
    .A2(_0525_),
    .B1(\bank_active[7] ),
    .Y(_0538_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(_0524_),
    .B(_0538_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand2_1 _1248_ (.A(net32),
    .B(_0639_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _1249_ (.A(_0281_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand4b_4 _1250_ (.A_N(_0323_),
    .B(_0420_),
    .C(_0540_),
    .D(_0067_),
    .Y(_0541_));
 sky130_fd_sc_hd__mux2i_2 _1251_ (.A0(\init_state[1] ),
    .A1(_0142_),
    .S(_0281_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(net118),
    .B(_0541_),
    .Y(_0543_));
 sky130_fd_sc_hd__o21ai_0 _1253_ (.A1(_0541_),
    .A2(_0542_),
    .B1(_0543_),
    .Y(_0040_));
 sky130_fd_sc_hd__nor2_1 _1254_ (.A(_0281_),
    .B(_0308_),
    .Y(_0544_));
 sky130_fd_sc_hd__a211oi_1 _1255_ (.A1(_0281_),
    .A2(_0121_),
    .B1(_0541_),
    .C1(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0619_),
    .A2(_0541_),
    .B1(_0545_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(net120),
    .B(_0541_),
    .Y(_0546_));
 sky130_fd_sc_hd__o31ai_1 _1258_ (.A1(_0298_),
    .A2(_0104_),
    .A3(_0541_),
    .B1(_0546_),
    .Y(_0042_));
 sky130_fd_sc_hd__nand2_1 _1259_ (.A(_0290_),
    .B(\burst_counter[0] ),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_0 _1260_ (.A1(_0290_),
    .A2(net28),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _1261_ (.A(_0050_),
    .B(_0377_),
    .Y(_0549_));
 sky130_fd_sc_hd__a22oi_1 _1262_ (.A1(_0313_),
    .A2(_0488_),
    .B1(_0549_),
    .B2(_0066_),
    .Y(_0550_));
 sky130_fd_sc_hd__and2_0 _1263_ (.A(_0152_),
    .B(_0153_),
    .X(_0551_));
 sky130_fd_sc_hd__a211o_1 _1264_ (.A1(_0164_),
    .A2(_0246_),
    .B1(_0251_),
    .C1(_0228_),
    .X(_0552_));
 sky130_fd_sc_hd__a2111oi_1 _1265_ (.A1(net17),
    .A2(_0162_),
    .B1(_0218_),
    .C1(_0231_),
    .D1(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2b_1 _1266_ (.A(_0193_),
    .B_N(_0203_),
    .Y(_0554_));
 sky130_fd_sc_hd__nor3_1 _1267_ (.A(_0317_),
    .B(_0288_),
    .C(_0550_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand4_1 _1268_ (.A(_0551_),
    .B(_0553_),
    .C(_0554_),
    .D(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand3_1 _1269_ (.A(_0116_),
    .B(_0274_),
    .C(_0275_),
    .Y(_0557_));
 sky130_fd_sc_hd__o31ai_1 _1270_ (.A1(net7),
    .A2(_0137_),
    .A3(_0138_),
    .B1(_0260_),
    .Y(_0558_));
 sky130_fd_sc_hd__o2bb2ai_1 _1271_ (.A1_N(net7),
    .A2_N(_0137_),
    .B1(_0180_),
    .B2(_0182_),
    .Y(_0559_));
 sky130_fd_sc_hd__or4b_1 _1272_ (.A(_0173_),
    .B(_0558_),
    .C(_0559_),
    .D_N(_0262_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_1 _1273_ (.A(_0126_),
    .B(_0214_),
    .Y(_0561_));
 sky130_fd_sc_hd__or4_1 _1274_ (.A(_0243_),
    .B(_0557_),
    .C(_0560_),
    .D(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__o22a_1 _1275_ (.A1(_0664_),
    .A2(_0550_),
    .B1(_0556_),
    .B2(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_6 _1276_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(\burst_counter[0] ),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_0 _1278_ (.A1(_0548_),
    .A2(_0564_),
    .B1(_0565_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _1279_ (.A(_0085_),
    .B(_0636_),
    .Y(_0566_));
 sky130_fd_sc_hd__o21ai_0 _1280_ (.A1(_0085_),
    .A2(net29),
    .B1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _1281_ (.A(\burst_counter[1] ),
    .B(_0564_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_0 _1282_ (.A1(_0564_),
    .A2(_0567_),
    .B1(_0568_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _1283_ (.A(\burst_counter[2] ),
    .B(_0564_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _1284_ (.A(_0084_),
    .B(_0637_),
    .Y(_0570_));
 sky130_fd_sc_hd__or3_1 _1285_ (.A(\burst_counter[2] ),
    .B(_0564_),
    .C(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__or3b_1 _1286_ (.A(_0564_),
    .B(_0084_),
    .C_N(net30),
    .X(_0572_));
 sky130_fd_sc_hd__nand3b_1 _1287_ (.A_N(_0637_),
    .B(\burst_counter[2] ),
    .C(_0085_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand4_1 _1288_ (.A(_0569_),
    .B(_0571_),
    .C(_0572_),
    .D(_0573_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2b_1 _1289_ (.A_N(_0290_),
    .B(net31),
    .Y(_0574_));
 sky130_fd_sc_hd__or3_1 _1290_ (.A(\burst_counter[2] ),
    .B(\burst_counter[1] ),
    .C(\burst_counter[0] ),
    .X(_0575_));
 sky130_fd_sc_hd__nand3_1 _1291_ (.A(_0085_),
    .B(\burst_counter[3] ),
    .C(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nor3b_1 _1292_ (.A(\burst_counter[3] ),
    .B(_0575_),
    .C_N(_0084_),
    .Y(_0577_));
 sky130_fd_sc_hd__mux2i_1 _1293_ (.A0(_0577_),
    .A1(\burst_counter[3] ),
    .S(_0564_),
    .Y(_0578_));
 sky130_fd_sc_hd__o211ai_1 _1294_ (.A1(_0564_),
    .A2(_0574_),
    .B1(_0576_),
    .C1(_0578_),
    .Y(_0046_));
 sky130_fd_sc_hd__nor2_1 _1295_ (.A(_0324_),
    .B(_0459_),
    .Y(_0579_));
 sky130_fd_sc_hd__o2111ai_1 _1296_ (.A1(_0298_),
    .A2(_0319_),
    .B1(_0579_),
    .C1(_0661_),
    .D1(_0300_),
    .Y(_0580_));
 sky130_fd_sc_hd__o21a_1 _1297_ (.A1(net199),
    .A2(_0579_),
    .B1(_0580_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0661_),
    .B(_0579_),
    .Y(_0581_));
 sky130_fd_sc_hd__o21ai_0 _1299_ (.A1(_0659_),
    .A2(_0579_),
    .B1(_0581_),
    .Y(_0048_));
 sky130_fd_sc_hd__a21o_1 _1300_ (.A1(\init_state[7] ),
    .A2(_0059_),
    .B1(net103),
    .X(_0049_));
 sky130_fd_sc_hd__nor2_1 _1301_ (.A(_0648_),
    .B(_0289_),
    .Y(net102));
 sky130_fd_sc_hd__inv_1 _1302_ (.A(cmd_reg_valid),
    .Y(net122));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(\init_state[7] ),
    .B(\init_state[3] ),
    .Y(_0582_));
 sky130_fd_sc_hd__a21boi_0 _1304_ (.A1(_0367_),
    .A2(_0582_),
    .B1_N(net36),
    .Y(net132));
 sky130_fd_sc_hd__ha_1 _1305_ (.A(_0618_),
    .B(_0619_),
    .COUT(_0620_),
    .SUM(_0621_));
 sky130_fd_sc_hd__ha_1 _1306_ (.A(_0618_),
    .B(net119),
    .COUT(_0622_),
    .SUM(_0623_));
 sky130_fd_sc_hd__ha_1 _1307_ (.A(net118),
    .B(_0619_),
    .COUT(_0624_),
    .SUM(_0625_));
 sky130_fd_sc_hd__ha_1 _1308_ (.A(net118),
    .B(net119),
    .COUT(_0626_),
    .SUM(_0627_));
 sky130_fd_sc_hd__ha_1 _1309_ (.A(_0628_),
    .B(_0620_),
    .COUT(_0629_),
    .SUM(_0630_));
 sky130_fd_sc_hd__ha_1 _1310_ (.A(net120),
    .B(_0620_),
    .COUT(_0631_),
    .SUM(_0632_));
 sky130_fd_sc_hd__ha_1 _1311_ (.A(_0633_),
    .B(_0634_),
    .COUT(_0635_),
    .SUM(_0636_));
 sky130_fd_sc_hd__ha_1 _1312_ (.A(_0633_),
    .B(_0634_),
    .COUT(_0637_),
    .SUM(_0638_));
 sky130_fd_sc_hd__ha_1 _1313_ (.A(_0639_),
    .B(_0640_),
    .COUT(_0641_),
    .SUM(_0642_));
 sky130_fd_sc_hd__ha_1 _1314_ (.A(_0640_),
    .B(\refresh_counter[1] ),
    .COUT(_0643_),
    .SUM(_0644_));
 sky130_fd_sc_hd__ha_1 _1315_ (.A(\refresh_counter[0] ),
    .B(\refresh_counter[1] ),
    .COUT(_0645_),
    .SUM(_0646_));
 sky130_fd_sc_hd__ha_1 _1316_ (.A(_0647_),
    .B(_0648_),
    .COUT(_0649_),
    .SUM(_0650_));
 sky130_fd_sc_hd__ha_1 _1317_ (.A(\timer[0] ),
    .B(_0648_),
    .COUT(_0651_),
    .SUM(_0652_));
 sky130_fd_sc_hd__ha_1 _1318_ (.A(_0647_),
    .B(_0653_),
    .COUT(_0654_),
    .SUM(_0655_));
 sky130_fd_sc_hd__ha_1 _1319_ (.A(\timer[0] ),
    .B(_0653_),
    .COUT(_0656_),
    .SUM(_0657_));
 sky130_fd_sc_hd__ha_1 _1320_ (.A(_0658_),
    .B(_0659_),
    .COUT(_0660_),
    .SUM(_0661_));
 sky130_fd_sc_hd__ha_1 _1321_ (.A(_0658_),
    .B(net200),
    .COUT(_0662_),
    .SUM(_0663_));
 sky130_fd_sc_hd__ha_2 _1322_ (.A(net199),
    .B(_0659_),
    .COUT(_0664_),
    .SUM(_0665_));
 sky130_fd_sc_hd__ha_1 _1323_ (.A(net199),
    .B(net200),
    .COUT(_0666_),
    .SUM(_0667_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__conb_1 _1328__211 (.HI(net212));
 sky130_fd_sc_hd__buf_4 _1326_ (.A(net202),
    .X(phy_bank_group[0]));
 sky130_fd_sc_hd__buf_4 _1327_ (.A(net203),
    .X(phy_bank_group[1]));
 sky130_fd_sc_hd__buf_4 _1328_ (.A(net212),
    .X(phy_cke));
 sky130_fd_sc_hd__clkbuf_1 _1329_ (.A(wr_mask[0]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 _1330_ (.A(wr_mask[1]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _1331_ (.A(wr_mask[2]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _1332_ (.A(wr_mask[3]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _1333_ (.A(wr_mask[4]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _1334_ (.A(wr_mask[5]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _1335_ (.A(wr_mask[6]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _1336_ (.A(wr_mask[7]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _1337_ (.A(net37),
    .X(phy_dq[0]));
 sky130_fd_sc_hd__clkbuf_1 _1338_ (.A(net48),
    .X(phy_dq[1]));
 sky130_fd_sc_hd__clkbuf_1 _1339_ (.A(net59),
    .X(phy_dq[2]));
 sky130_fd_sc_hd__clkbuf_1 _1340_ (.A(net70),
    .X(phy_dq[3]));
 sky130_fd_sc_hd__clkbuf_1 _1341_ (.A(net81),
    .X(phy_dq[4]));
 sky130_fd_sc_hd__clkbuf_1 _1342_ (.A(net92),
    .X(phy_dq[5]));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(net97),
    .X(phy_dq[6]));
 sky130_fd_sc_hd__clkbuf_1 _1344_ (.A(net98),
    .X(phy_dq[7]));
 sky130_fd_sc_hd__clkbuf_1 _1345_ (.A(net99),
    .X(phy_dq[8]));
 sky130_fd_sc_hd__clkbuf_1 _1346_ (.A(net100),
    .X(phy_dq[9]));
 sky130_fd_sc_hd__clkbuf_1 _1347_ (.A(net38),
    .X(phy_dq[10]));
 sky130_fd_sc_hd__clkbuf_1 _1348_ (.A(net39),
    .X(phy_dq[11]));
 sky130_fd_sc_hd__clkbuf_1 _1349_ (.A(net40),
    .X(phy_dq[12]));
 sky130_fd_sc_hd__clkbuf_1 _1350_ (.A(net41),
    .X(phy_dq[13]));
 sky130_fd_sc_hd__clkbuf_1 _1351_ (.A(net42),
    .X(phy_dq[14]));
 sky130_fd_sc_hd__clkbuf_1 _1352_ (.A(net43),
    .X(phy_dq[15]));
 sky130_fd_sc_hd__clkbuf_1 _1353_ (.A(net44),
    .X(phy_dq[16]));
 sky130_fd_sc_hd__clkbuf_1 _1354_ (.A(net45),
    .X(phy_dq[17]));
 sky130_fd_sc_hd__clkbuf_1 _1355_ (.A(net46),
    .X(phy_dq[18]));
 sky130_fd_sc_hd__clkbuf_1 _1356_ (.A(net47),
    .X(phy_dq[19]));
 sky130_fd_sc_hd__clkbuf_1 _1357_ (.A(net49),
    .X(phy_dq[20]));
 sky130_fd_sc_hd__clkbuf_1 _1358_ (.A(net50),
    .X(phy_dq[21]));
 sky130_fd_sc_hd__clkbuf_1 _1359_ (.A(net51),
    .X(phy_dq[22]));
 sky130_fd_sc_hd__clkbuf_1 _1360_ (.A(net52),
    .X(phy_dq[23]));
 sky130_fd_sc_hd__clkbuf_1 _1361_ (.A(net53),
    .X(phy_dq[24]));
 sky130_fd_sc_hd__clkbuf_1 _1362_ (.A(net54),
    .X(phy_dq[25]));
 sky130_fd_sc_hd__clkbuf_1 _1363_ (.A(net55),
    .X(phy_dq[26]));
 sky130_fd_sc_hd__clkbuf_1 _1364_ (.A(net56),
    .X(phy_dq[27]));
 sky130_fd_sc_hd__clkbuf_1 _1365_ (.A(net57),
    .X(phy_dq[28]));
 sky130_fd_sc_hd__clkbuf_1 _1366_ (.A(net58),
    .X(phy_dq[29]));
 sky130_fd_sc_hd__clkbuf_1 _1367_ (.A(net60),
    .X(phy_dq[30]));
 sky130_fd_sc_hd__clkbuf_1 _1368_ (.A(net61),
    .X(phy_dq[31]));
 sky130_fd_sc_hd__clkbuf_1 _1369_ (.A(net62),
    .X(phy_dq[32]));
 sky130_fd_sc_hd__clkbuf_1 _1370_ (.A(net63),
    .X(phy_dq[33]));
 sky130_fd_sc_hd__clkbuf_1 _1371_ (.A(net64),
    .X(phy_dq[34]));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(net65),
    .X(phy_dq[35]));
 sky130_fd_sc_hd__clkbuf_1 _1373_ (.A(net66),
    .X(phy_dq[36]));
 sky130_fd_sc_hd__clkbuf_1 _1374_ (.A(net67),
    .X(phy_dq[37]));
 sky130_fd_sc_hd__clkbuf_1 _1375_ (.A(net68),
    .X(phy_dq[38]));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(net69),
    .X(phy_dq[39]));
 sky130_fd_sc_hd__clkbuf_1 _1377_ (.A(net71),
    .X(phy_dq[40]));
 sky130_fd_sc_hd__clkbuf_1 _1378_ (.A(net72),
    .X(phy_dq[41]));
 sky130_fd_sc_hd__clkbuf_1 _1379_ (.A(net73),
    .X(phy_dq[42]));
 sky130_fd_sc_hd__clkbuf_1 _1380_ (.A(net74),
    .X(phy_dq[43]));
 sky130_fd_sc_hd__clkbuf_1 _1381_ (.A(net75),
    .X(phy_dq[44]));
 sky130_fd_sc_hd__clkbuf_1 _1382_ (.A(net76),
    .X(phy_dq[45]));
 sky130_fd_sc_hd__clkbuf_1 _1383_ (.A(net77),
    .X(phy_dq[46]));
 sky130_fd_sc_hd__clkbuf_1 _1384_ (.A(net78),
    .X(phy_dq[47]));
 sky130_fd_sc_hd__clkbuf_1 _1385_ (.A(net79),
    .X(phy_dq[48]));
 sky130_fd_sc_hd__clkbuf_1 _1386_ (.A(net80),
    .X(phy_dq[49]));
 sky130_fd_sc_hd__clkbuf_1 _1387_ (.A(net82),
    .X(phy_dq[50]));
 sky130_fd_sc_hd__clkbuf_1 _1388_ (.A(net83),
    .X(phy_dq[51]));
 sky130_fd_sc_hd__clkbuf_1 _1389_ (.A(net84),
    .X(phy_dq[52]));
 sky130_fd_sc_hd__clkbuf_1 _1390_ (.A(net85),
    .X(phy_dq[53]));
 sky130_fd_sc_hd__clkbuf_1 _1391_ (.A(net86),
    .X(phy_dq[54]));
 sky130_fd_sc_hd__clkbuf_1 _1392_ (.A(net87),
    .X(phy_dq[55]));
 sky130_fd_sc_hd__clkbuf_1 _1393_ (.A(net88),
    .X(phy_dq[56]));
 sky130_fd_sc_hd__clkbuf_1 _1394_ (.A(net89),
    .X(phy_dq[57]));
 sky130_fd_sc_hd__clkbuf_1 _1395_ (.A(net90),
    .X(phy_dq[58]));
 sky130_fd_sc_hd__clkbuf_1 _1396_ (.A(net91),
    .X(phy_dq[59]));
 sky130_fd_sc_hd__clkbuf_1 _1397_ (.A(net93),
    .X(phy_dq[60]));
 sky130_fd_sc_hd__clkbuf_1 _1398_ (.A(net94),
    .X(phy_dq[61]));
 sky130_fd_sc_hd__clkbuf_1 _1399_ (.A(net95),
    .X(phy_dq[62]));
 sky130_fd_sc_hd__clkbuf_1 _1400_ (.A(net96),
    .X(phy_dq[63]));
 sky130_fd_sc_hd__buf_4 _1401_ (.A(net204),
    .X(phy_dqs_n[0]));
 sky130_fd_sc_hd__buf_4 _1402_ (.A(net205),
    .X(phy_dqs_n[1]));
 sky130_fd_sc_hd__buf_4 _1403_ (.A(net206),
    .X(phy_dqs_n[2]));
 sky130_fd_sc_hd__buf_4 _1404_ (.A(net207),
    .X(phy_dqs_n[3]));
 sky130_fd_sc_hd__buf_4 _1405_ (.A(net208),
    .X(phy_dqs_n[4]));
 sky130_fd_sc_hd__buf_4 _1406_ (.A(net209),
    .X(phy_dqs_n[5]));
 sky130_fd_sc_hd__buf_4 _1407_ (.A(net210),
    .X(phy_dqs_n[6]));
 sky130_fd_sc_hd__buf_4 _1408_ (.A(net211),
    .X(phy_dqs_n[7]));
 sky130_fd_sc_hd__buf_4 _1409_ (.A(net213),
    .X(phy_dqs_p[0]));
 sky130_fd_sc_hd__buf_4 _1410_ (.A(net214),
    .X(phy_dqs_p[1]));
 sky130_fd_sc_hd__buf_4 _1411_ (.A(net215),
    .X(phy_dqs_p[2]));
 sky130_fd_sc_hd__buf_4 _1412_ (.A(net216),
    .X(phy_dqs_p[3]));
 sky130_fd_sc_hd__buf_4 _1413_ (.A(net217),
    .X(phy_dqs_p[4]));
 sky130_fd_sc_hd__buf_4 _1414_ (.A(net218),
    .X(phy_dqs_p[5]));
 sky130_fd_sc_hd__buf_4 _1415_ (.A(net219),
    .X(phy_dqs_p[6]));
 sky130_fd_sc_hd__buf_4 _1416_ (.A(net220),
    .X(phy_dqs_p[7]));
 sky130_fd_sc_hd__buf_4 _1417_ (.A(net221),
    .X(phy_odt));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][0]$_DFFE_PP_  (.D(net104),
    .DE(_0016_),
    .Q(\active_row[0][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][10]$_DFFE_PP_  (.D(net105),
    .DE(_0016_),
    .Q(\active_row[0][10] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][11]$_DFFE_PP_  (.D(net106),
    .DE(_0016_),
    .Q(\active_row[0][11] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][12]$_DFFE_PP_  (.D(net107),
    .DE(_0016_),
    .Q(\active_row[0][12] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][13]$_DFFE_PP_  (.D(net108),
    .DE(_0016_),
    .Q(\active_row[0][13] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][1]$_DFFE_PP_  (.D(net109),
    .DE(_0016_),
    .Q(\active_row[0][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][2]$_DFFE_PP_  (.D(net110),
    .DE(_0016_),
    .Q(\active_row[0][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][3]$_DFFE_PP_  (.D(net111),
    .DE(_0016_),
    .Q(\active_row[0][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][4]$_DFFE_PP_  (.D(net112),
    .DE(_0016_),
    .Q(\active_row[0][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][5]$_DFFE_PP_  (.D(net113),
    .DE(_0016_),
    .Q(\active_row[0][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][6]$_DFFE_PP_  (.D(net114),
    .DE(_0016_),
    .Q(\active_row[0][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][7]$_DFFE_PP_  (.D(net115),
    .DE(_0016_),
    .Q(\active_row[0][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][8]$_DFFE_PP_  (.D(net116),
    .DE(_0016_),
    .Q(\active_row[0][8] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[0][9]$_DFFE_PP_  (.D(net117),
    .DE(_0016_),
    .Q(\active_row[0][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][0]$_DFFE_PP_  (.D(net104),
    .DE(_0015_),
    .Q(\active_row[1][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][10]$_DFFE_PP_  (.D(net105),
    .DE(_0015_),
    .Q(\active_row[1][10] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][11]$_DFFE_PP_  (.D(net106),
    .DE(_0015_),
    .Q(\active_row[1][11] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][12]$_DFFE_PP_  (.D(net107),
    .DE(_0015_),
    .Q(\active_row[1][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][13]$_DFFE_PP_  (.D(net108),
    .DE(_0015_),
    .Q(\active_row[1][13] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][1]$_DFFE_PP_  (.D(net109),
    .DE(_0015_),
    .Q(\active_row[1][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][2]$_DFFE_PP_  (.D(net110),
    .DE(_0015_),
    .Q(\active_row[1][2] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][3]$_DFFE_PP_  (.D(net111),
    .DE(_0015_),
    .Q(\active_row[1][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][4]$_DFFE_PP_  (.D(net112),
    .DE(_0015_),
    .Q(\active_row[1][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][5]$_DFFE_PP_  (.D(net113),
    .DE(_0015_),
    .Q(\active_row[1][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][6]$_DFFE_PP_  (.D(net114),
    .DE(_0015_),
    .Q(\active_row[1][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][7]$_DFFE_PP_  (.D(net115),
    .DE(_0015_),
    .Q(\active_row[1][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][8]$_DFFE_PP_  (.D(net116),
    .DE(_0015_),
    .Q(\active_row[1][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[1][9]$_DFFE_PP_  (.D(net117),
    .DE(_0015_),
    .Q(\active_row[1][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][0]$_DFFE_PP_  (.D(net104),
    .DE(_0014_),
    .Q(\active_row[2][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][10]$_DFFE_PP_  (.D(net105),
    .DE(_0014_),
    .Q(\active_row[2][10] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][11]$_DFFE_PP_  (.D(net106),
    .DE(_0014_),
    .Q(\active_row[2][11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][12]$_DFFE_PP_  (.D(net107),
    .DE(_0014_),
    .Q(\active_row[2][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][13]$_DFFE_PP_  (.D(net108),
    .DE(_0014_),
    .Q(\active_row[2][13] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][1]$_DFFE_PP_  (.D(net109),
    .DE(_0014_),
    .Q(\active_row[2][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][2]$_DFFE_PP_  (.D(net110),
    .DE(_0014_),
    .Q(\active_row[2][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][3]$_DFFE_PP_  (.D(net111),
    .DE(_0014_),
    .Q(\active_row[2][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][4]$_DFFE_PP_  (.D(net112),
    .DE(_0014_),
    .Q(\active_row[2][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][5]$_DFFE_PP_  (.D(net113),
    .DE(_0014_),
    .Q(\active_row[2][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][6]$_DFFE_PP_  (.D(net114),
    .DE(_0014_),
    .Q(\active_row[2][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][7]$_DFFE_PP_  (.D(net115),
    .DE(_0014_),
    .Q(\active_row[2][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][8]$_DFFE_PP_  (.D(net116),
    .DE(_0014_),
    .Q(\active_row[2][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[2][9]$_DFFE_PP_  (.D(net117),
    .DE(_0014_),
    .Q(\active_row[2][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][0]$_DFFE_PP_  (.D(net104),
    .DE(_0013_),
    .Q(\active_row[3][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][10]$_DFFE_PP_  (.D(net105),
    .DE(_0013_),
    .Q(\active_row[3][10] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][11]$_DFFE_PP_  (.D(net106),
    .DE(_0013_),
    .Q(\active_row[3][11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][12]$_DFFE_PP_  (.D(net107),
    .DE(_0013_),
    .Q(\active_row[3][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][13]$_DFFE_PP_  (.D(net108),
    .DE(_0013_),
    .Q(\active_row[3][13] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][1]$_DFFE_PP_  (.D(net109),
    .DE(_0013_),
    .Q(\active_row[3][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][2]$_DFFE_PP_  (.D(net110),
    .DE(_0013_),
    .Q(\active_row[3][2] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][3]$_DFFE_PP_  (.D(net111),
    .DE(_0013_),
    .Q(\active_row[3][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][4]$_DFFE_PP_  (.D(net112),
    .DE(_0013_),
    .Q(\active_row[3][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][5]$_DFFE_PP_  (.D(net113),
    .DE(_0013_),
    .Q(\active_row[3][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][6]$_DFFE_PP_  (.D(net114),
    .DE(_0013_),
    .Q(\active_row[3][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][7]$_DFFE_PP_  (.D(net115),
    .DE(_0013_),
    .Q(\active_row[3][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][8]$_DFFE_PP_  (.D(net116),
    .DE(_0013_),
    .Q(\active_row[3][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[3][9]$_DFFE_PP_  (.D(net117),
    .DE(_0013_),
    .Q(\active_row[3][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][0]$_DFFE_PP_  (.D(net104),
    .DE(_0012_),
    .Q(\active_row[4][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][10]$_DFFE_PP_  (.D(net105),
    .DE(_0012_),
    .Q(\active_row[4][10] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][11]$_DFFE_PP_  (.D(net106),
    .DE(_0012_),
    .Q(\active_row[4][11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][12]$_DFFE_PP_  (.D(net107),
    .DE(_0012_),
    .Q(\active_row[4][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][13]$_DFFE_PP_  (.D(net108),
    .DE(_0012_),
    .Q(\active_row[4][13] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][1]$_DFFE_PP_  (.D(net109),
    .DE(_0012_),
    .Q(\active_row[4][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][2]$_DFFE_PP_  (.D(net110),
    .DE(_0012_),
    .Q(\active_row[4][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][3]$_DFFE_PP_  (.D(net111),
    .DE(_0012_),
    .Q(\active_row[4][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][4]$_DFFE_PP_  (.D(net112),
    .DE(_0012_),
    .Q(\active_row[4][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][5]$_DFFE_PP_  (.D(net113),
    .DE(_0012_),
    .Q(\active_row[4][5] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][6]$_DFFE_PP_  (.D(net114),
    .DE(_0012_),
    .Q(\active_row[4][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][7]$_DFFE_PP_  (.D(net115),
    .DE(_0012_),
    .Q(\active_row[4][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][8]$_DFFE_PP_  (.D(net116),
    .DE(_0012_),
    .Q(\active_row[4][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[4][9]$_DFFE_PP_  (.D(net117),
    .DE(_0012_),
    .Q(\active_row[4][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][0]$_DFFE_PP_  (.D(net104),
    .DE(_0011_),
    .Q(\active_row[5][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][10]$_DFFE_PP_  (.D(net105),
    .DE(_0011_),
    .Q(\active_row[5][10] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][11]$_DFFE_PP_  (.D(net106),
    .DE(_0011_),
    .Q(\active_row[5][11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][12]$_DFFE_PP_  (.D(net107),
    .DE(_0011_),
    .Q(\active_row[5][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][13]$_DFFE_PP_  (.D(net108),
    .DE(_0011_),
    .Q(\active_row[5][13] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][1]$_DFFE_PP_  (.D(net109),
    .DE(_0011_),
    .Q(\active_row[5][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][2]$_DFFE_PP_  (.D(net110),
    .DE(_0011_),
    .Q(\active_row[5][2] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][3]$_DFFE_PP_  (.D(net111),
    .DE(_0011_),
    .Q(\active_row[5][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][4]$_DFFE_PP_  (.D(net112),
    .DE(_0011_),
    .Q(\active_row[5][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][5]$_DFFE_PP_  (.D(net113),
    .DE(_0011_),
    .Q(\active_row[5][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][6]$_DFFE_PP_  (.D(net114),
    .DE(_0011_),
    .Q(\active_row[5][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][7]$_DFFE_PP_  (.D(net115),
    .DE(_0011_),
    .Q(\active_row[5][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][8]$_DFFE_PP_  (.D(net116),
    .DE(_0011_),
    .Q(\active_row[5][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[5][9]$_DFFE_PP_  (.D(net117),
    .DE(_0011_),
    .Q(\active_row[5][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][0]$_DFFE_PP_  (.D(net104),
    .DE(_0010_),
    .Q(\active_row[6][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][10]$_DFFE_PP_  (.D(net105),
    .DE(_0010_),
    .Q(\active_row[6][10] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][11]$_DFFE_PP_  (.D(net106),
    .DE(_0010_),
    .Q(\active_row[6][11] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][12]$_DFFE_PP_  (.D(net107),
    .DE(_0010_),
    .Q(\active_row[6][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][13]$_DFFE_PP_  (.D(net108),
    .DE(_0010_),
    .Q(\active_row[6][13] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][1]$_DFFE_PP_  (.D(net109),
    .DE(_0010_),
    .Q(\active_row[6][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][2]$_DFFE_PP_  (.D(net110),
    .DE(_0010_),
    .Q(\active_row[6][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][3]$_DFFE_PP_  (.D(net111),
    .DE(_0010_),
    .Q(\active_row[6][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][4]$_DFFE_PP_  (.D(net112),
    .DE(_0010_),
    .Q(\active_row[6][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][5]$_DFFE_PP_  (.D(net113),
    .DE(_0010_),
    .Q(\active_row[6][5] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][6]$_DFFE_PP_  (.D(net114),
    .DE(_0010_),
    .Q(\active_row[6][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][7]$_DFFE_PP_  (.D(net115),
    .DE(_0010_),
    .Q(\active_row[6][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][8]$_DFFE_PP_  (.D(net116),
    .DE(_0010_),
    .Q(\active_row[6][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[6][9]$_DFFE_PP_  (.D(net117),
    .DE(_0010_),
    .Q(\active_row[6][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][0]$_DFFE_PP_  (.D(net104),
    .DE(_0009_),
    .Q(\active_row[7][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][10]$_DFFE_PP_  (.D(net105),
    .DE(_0009_),
    .Q(\active_row[7][10] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][11]$_DFFE_PP_  (.D(net106),
    .DE(_0009_),
    .Q(\active_row[7][11] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][12]$_DFFE_PP_  (.D(net107),
    .DE(_0009_),
    .Q(\active_row[7][12] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][13]$_DFFE_PP_  (.D(net108),
    .DE(_0009_),
    .Q(\active_row[7][13] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][1]$_DFFE_PP_  (.D(net109),
    .DE(_0009_),
    .Q(\active_row[7][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][2]$_DFFE_PP_  (.D(net110),
    .DE(_0009_),
    .Q(\active_row[7][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][3]$_DFFE_PP_  (.D(net111),
    .DE(_0009_),
    .Q(\active_row[7][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][4]$_DFFE_PP_  (.D(net112),
    .DE(_0009_),
    .Q(\active_row[7][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][5]$_DFFE_PP_  (.D(net113),
    .DE(_0009_),
    .Q(\active_row[7][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][6]$_DFFE_PP_  (.D(net114),
    .DE(_0009_),
    .Q(\active_row[7][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][7]$_DFFE_PP_  (.D(net115),
    .DE(_0009_),
    .Q(\active_row[7][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][8]$_DFFE_PP_  (.D(net116),
    .DE(_0009_),
    .Q(\active_row[7][8] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \active_row[7][9]$_DFFE_PP_  (.D(net117),
    .DE(_0009_),
    .Q(\active_row[7][9] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[0]$_DFFE_PN0P_  (.D(_0018_),
    .Q(net104),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[10]$_DFFE_PN0P_  (.D(_0019_),
    .Q(net105),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[11]$_DFFE_PN0P_  (.D(_0020_),
    .Q(net106),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[12]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net107),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[13]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net108),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[1]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net109),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[2]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net110),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[3]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net111),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[4]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net112),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[5]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net113),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[6]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net114),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[7]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net115),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[8]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net116),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_reg[9]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net117),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[0]$_DFFE_PN0P_  (.D(_0032_),
    .Q(\bank_active[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[1]$_DFFE_PN0P_  (.D(_0033_),
    .Q(\bank_active[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[2]$_DFFE_PN0P_  (.D(_0034_),
    .Q(\bank_active[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[3]$_DFFE_PN0P_  (.D(_0035_),
    .Q(\bank_active[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[4]$_DFFE_PN0P_  (.D(_0036_),
    .Q(\bank_active[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[5]$_DFFE_PN0P_  (.D(_0037_),
    .Q(\bank_active[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[6]$_DFFE_PN0P_  (.D(_0038_),
    .Q(\bank_active[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \bank_active[7]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\bank_active[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \bank_reg[0]$_DFFE_PN0P_  (.D(_0040_),
    .Q(net118),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \bank_reg[1]$_DFFE_PN0P_  (.D(_0041_),
    .Q(net119),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \bank_reg[2]$_DFFE_PN0P_  (.D(_0042_),
    .Q(net120),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \burst_counter[0]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\burst_counter[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \burst_counter[1]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\burst_counter[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \burst_counter[2]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\burst_counter[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \burst_counter[3]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\burst_counter[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfstp_1 \cmd_reg[0]$_DFF_PN1_  (.D(_0583_),
    .Q(net133),
    .SET_B(net36),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfstp_1 \cmd_reg[1]$_DFF_PN1_  (.D(_0584_),
    .Q(net121),
    .SET_B(net36),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfstp_1 \cmd_reg[2]$_DFF_PN1_  (.D(_0585_),
    .Q(net131),
    .SET_B(net36),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \cmd_reg_valid$_DFF_PN0_  (.D(net222),
    .Q(cmd_reg_valid),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \curr_state[0]$_DFFE_PN0P_  (.D(_0047_),
    .Q(net199),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \curr_state[1]$_DFFE_PN0P_  (.D(_0048_),
    .Q(net200),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_done_reg$_DFFE_PN0P_  (.D(_0049_),
    .Q(net103),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfstp_1 \init_state[0]$_DFF_PN1_  (.D(_0001_),
    .Q(\init_state[0] ),
    .SET_B(net36),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \init_state[1]$_DFF_PN0_  (.D(_0002_),
    .Q(\init_state[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_state[2]$_DFF_PN0_  (.D(_0003_),
    .Q(\init_state[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_state[3]$_DFF_PN0_  (.D(_0004_),
    .Q(\init_state[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_state[4]$_DFF_PN0_  (.D(_0005_),
    .Q(\init_state[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_state[5]$_DFF_PN0_  (.D(_0006_),
    .Q(\init_state[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \init_state[6]$_DFF_PN0_  (.D(_0007_),
    .Q(\init_state[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \init_state[7]$_DFF_PN0_  (.D(_0008_),
    .Q(\init_state[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[0]$_DFFE_PP_  (.D(net37),
    .DE(_0017_),
    .Q(net134),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[10]$_DFFE_PP_  (.D(net38),
    .DE(_0017_),
    .Q(net135),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[11]$_DFFE_PP_  (.D(net39),
    .DE(_0017_),
    .Q(net136),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[12]$_DFFE_PP_  (.D(net40),
    .DE(_0017_),
    .Q(net137),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[13]$_DFFE_PP_  (.D(net41),
    .DE(_0017_),
    .Q(net138),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[14]$_DFFE_PP_  (.D(net42),
    .DE(_0017_),
    .Q(net139),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[15]$_DFFE_PP_  (.D(net43),
    .DE(_0017_),
    .Q(net140),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[16]$_DFFE_PP_  (.D(net44),
    .DE(_0017_),
    .Q(net141),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[17]$_DFFE_PP_  (.D(net45),
    .DE(_0017_),
    .Q(net142),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[18]$_DFFE_PP_  (.D(net46),
    .DE(_0017_),
    .Q(net143),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[19]$_DFFE_PP_  (.D(net47),
    .DE(_0017_),
    .Q(net144),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[1]$_DFFE_PP_  (.D(net48),
    .DE(_0017_),
    .Q(net145),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[20]$_DFFE_PP_  (.D(net49),
    .DE(_0017_),
    .Q(net146),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[21]$_DFFE_PP_  (.D(net50),
    .DE(_0017_),
    .Q(net147),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[22]$_DFFE_PP_  (.D(net51),
    .DE(_0017_),
    .Q(net148),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[23]$_DFFE_PP_  (.D(net52),
    .DE(_0017_),
    .Q(net149),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[24]$_DFFE_PP_  (.D(net53),
    .DE(_0017_),
    .Q(net150),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[25]$_DFFE_PP_  (.D(net54),
    .DE(_0017_),
    .Q(net151),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[26]$_DFFE_PP_  (.D(net55),
    .DE(_0017_),
    .Q(net152),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[27]$_DFFE_PP_  (.D(net56),
    .DE(_0017_),
    .Q(net153),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[28]$_DFFE_PP_  (.D(net57),
    .DE(_0017_),
    .Q(net154),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[29]$_DFFE_PP_  (.D(net58),
    .DE(_0017_),
    .Q(net155),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[2]$_DFFE_PP_  (.D(net59),
    .DE(_0017_),
    .Q(net156),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[30]$_DFFE_PP_  (.D(net60),
    .DE(_0017_),
    .Q(net157),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[31]$_DFFE_PP_  (.D(net61),
    .DE(_0017_),
    .Q(net158),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[32]$_DFFE_PP_  (.D(net62),
    .DE(_0017_),
    .Q(net159),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[33]$_DFFE_PP_  (.D(net63),
    .DE(_0017_),
    .Q(net160),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[34]$_DFFE_PP_  (.D(net64),
    .DE(_0017_),
    .Q(net161),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[35]$_DFFE_PP_  (.D(net65),
    .DE(_0017_),
    .Q(net162),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[36]$_DFFE_PP_  (.D(net66),
    .DE(_0017_),
    .Q(net163),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[37]$_DFFE_PP_  (.D(net67),
    .DE(_0017_),
    .Q(net164),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[38]$_DFFE_PP_  (.D(net68),
    .DE(_0017_),
    .Q(net165),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[39]$_DFFE_PP_  (.D(net69),
    .DE(_0017_),
    .Q(net166),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[3]$_DFFE_PP_  (.D(net70),
    .DE(_0017_),
    .Q(net167),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[40]$_DFFE_PP_  (.D(net71),
    .DE(_0017_),
    .Q(net168),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[41]$_DFFE_PP_  (.D(net72),
    .DE(_0017_),
    .Q(net169),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[42]$_DFFE_PP_  (.D(net73),
    .DE(_0017_),
    .Q(net170),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[43]$_DFFE_PP_  (.D(net74),
    .DE(_0017_),
    .Q(net171),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[44]$_DFFE_PP_  (.D(net75),
    .DE(_0017_),
    .Q(net172),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[45]$_DFFE_PP_  (.D(net76),
    .DE(_0017_),
    .Q(net173),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[46]$_DFFE_PP_  (.D(net77),
    .DE(_0017_),
    .Q(net174),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[47]$_DFFE_PP_  (.D(net78),
    .DE(_0017_),
    .Q(net175),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[48]$_DFFE_PP_  (.D(net79),
    .DE(_0017_),
    .Q(net176),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[49]$_DFFE_PP_  (.D(net80),
    .DE(_0017_),
    .Q(net177),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[4]$_DFFE_PP_  (.D(net81),
    .DE(_0017_),
    .Q(net178),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[50]$_DFFE_PP_  (.D(net82),
    .DE(_0017_),
    .Q(net179),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[51]$_DFFE_PP_  (.D(net83),
    .DE(_0017_),
    .Q(net180),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[52]$_DFFE_PP_  (.D(net84),
    .DE(_0017_),
    .Q(net181),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[53]$_DFFE_PP_  (.D(net85),
    .DE(_0017_),
    .Q(net182),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[54]$_DFFE_PP_  (.D(net86),
    .DE(_0017_),
    .Q(net183),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[55]$_DFFE_PP_  (.D(net87),
    .DE(_0017_),
    .Q(net184),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[56]$_DFFE_PP_  (.D(net88),
    .DE(_0017_),
    .Q(net185),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[57]$_DFFE_PP_  (.D(net89),
    .DE(_0017_),
    .Q(net186),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[58]$_DFFE_PP_  (.D(net90),
    .DE(_0017_),
    .Q(net187),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[59]$_DFFE_PP_  (.D(net91),
    .DE(_0017_),
    .Q(net188),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[5]$_DFFE_PP_  (.D(net92),
    .DE(_0017_),
    .Q(net189),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[60]$_DFFE_PP_  (.D(net93),
    .DE(_0017_),
    .Q(net190),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[61]$_DFFE_PP_  (.D(net94),
    .DE(_0017_),
    .Q(net191),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[62]$_DFFE_PP_  (.D(net95),
    .DE(_0017_),
    .Q(net192),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[63]$_DFFE_PP_  (.D(net96),
    .DE(_0017_),
    .Q(net193),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[6]$_DFFE_PP_  (.D(net97),
    .DE(_0017_),
    .Q(net194),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[7]$_DFFE_PP_  (.D(net98),
    .DE(_0017_),
    .Q(net195),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[8]$_DFFE_PP_  (.D(net99),
    .DE(_0017_),
    .Q(net196),
    .CLK(net34));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[9]$_DFFE_PP_  (.D(net100),
    .DE(_0017_),
    .Q(net197),
    .CLK(net34));
 sky130_fd_sc_hd__dfrtp_1 \rd_valid_reg$_DFF_PN0_  (.D(_0000_),
    .Q(net198),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[0]$_DFF_PN0_  (.D(_0586_),
    .Q(\refresh_counter[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[10]$_DFF_PN0_  (.D(_0587_),
    .Q(\refresh_counter[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[11]$_DFF_PN0_  (.D(_0588_),
    .Q(\refresh_counter[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[12]$_DFF_PN0_  (.D(_0589_),
    .Q(\refresh_counter[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[13]$_DFF_PN0_  (.D(_0590_),
    .Q(\refresh_counter[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[14]$_DFF_PN0_  (.D(_0591_),
    .Q(\refresh_counter[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[15]$_DFF_PN0_  (.D(_0592_),
    .Q(\refresh_counter[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[1]$_DFF_PN0_  (.D(_0593_),
    .Q(\refresh_counter[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[2]$_DFF_PN0_  (.D(_0594_),
    .Q(\refresh_counter[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[3]$_DFF_PN0_  (.D(_0595_),
    .Q(\refresh_counter[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[4]$_DFF_PN0_  (.D(_0596_),
    .Q(\refresh_counter[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[5]$_DFF_PN0_  (.D(_0597_),
    .Q(\refresh_counter[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[6]$_DFF_PN0_  (.D(_0598_),
    .Q(\refresh_counter[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[7]$_DFF_PN0_  (.D(_0599_),
    .Q(\refresh_counter[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[8]$_DFF_PN0_  (.D(_0600_),
    .Q(\refresh_counter[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \refresh_counter[9]$_DFF_PN0_  (.D(_0601_),
    .Q(\refresh_counter[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[0]$_DFF_PN0_  (.D(_0602_),
    .Q(\timer[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[10]$_DFF_PN0_  (.D(_0603_),
    .Q(\timer[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[11]$_DFF_PN0_  (.D(_0604_),
    .Q(\timer[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[12]$_DFF_PN0_  (.D(_0605_),
    .Q(\timer[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[13]$_DFF_PN0_  (.D(_0606_),
    .Q(\timer[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[14]$_DFF_PN0_  (.D(_0607_),
    .Q(\timer[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[15]$_DFF_PN0_  (.D(_0608_),
    .Q(\timer[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \timer[1]$_DFF_PN0_  (.D(_0609_),
    .Q(\timer[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[2]$_DFF_PN0_  (.D(_0610_),
    .Q(\timer[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[3]$_DFF_PN0_  (.D(_0611_),
    .Q(\timer[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[4]$_DFF_PN0_  (.D(_0612_),
    .Q(\timer[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[5]$_DFF_PN0_  (.D(_0613_),
    .Q(\timer[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[6]$_DFF_PN0_  (.D(_0614_),
    .Q(\timer[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[7]$_DFF_PN0_  (.D(_0615_),
    .Q(\timer[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[8]$_DFF_PN0_  (.D(_0616_),
    .Q(\timer[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \timer[9]$_DFF_PN0_  (.D(_0617_),
    .Q(\timer[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ready_reg$_DFF_PN0_  (.D(_0670_),
    .Q(net201),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net36),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_274 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(cmd_addr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(cmd_addr[11]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(cmd_addr[13]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(cmd_addr[14]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(cmd_addr[15]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input6 (.A(cmd_addr[16]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(cmd_addr[17]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(cmd_addr[18]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(cmd_addr[19]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(cmd_addr[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(cmd_addr[20]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(cmd_addr[21]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(cmd_addr[22]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(cmd_addr[23]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(cmd_addr[24]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(cmd_addr[25]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(cmd_addr[26]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(cmd_addr[27]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(cmd_addr[2]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(cmd_addr[3]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(cmd_addr[4]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(cmd_addr[5]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(cmd_addr[6]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(cmd_addr[7]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(cmd_addr[8]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(cmd_addr[9]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(cmd_burst_len[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(cmd_burst_len[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(cmd_burst_len[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(cmd_burst_len[3]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(cmd_valid),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(cmd_write),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input33 (.A(phy_clk),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(rd_ready),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(net223),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(wr_data[0]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(wr_data[10]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(wr_data[11]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(wr_data[12]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(wr_data[13]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(wr_data[14]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(wr_data[15]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(wr_data[16]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(wr_data[17]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(wr_data[18]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(wr_data[19]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(wr_data[1]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(wr_data[20]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(wr_data[21]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(wr_data[22]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(wr_data[23]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(wr_data[24]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(wr_data[25]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(wr_data[26]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(wr_data[27]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(wr_data[28]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(wr_data[29]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(wr_data[2]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(wr_data[30]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(wr_data[31]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(wr_data[32]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(wr_data[33]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(wr_data[34]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(wr_data[35]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(wr_data[36]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wr_data[37]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wr_data[38]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(wr_data[39]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(wr_data[3]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(wr_data[40]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(wr_data[41]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(wr_data[42]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(wr_data[43]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(wr_data[44]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(wr_data[45]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(wr_data[46]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(wr_data[47]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(wr_data[48]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(wr_data[49]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(wr_data[4]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(wr_data[50]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(wr_data[51]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(wr_data[52]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(wr_data[53]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(wr_data[54]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(wr_data[55]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(wr_data[56]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(wr_data[57]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(wr_data[58]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(wr_data[59]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(wr_data[5]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(wr_data[60]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(wr_data[61]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(wr_data[62]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(wr_data[63]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(wr_data[6]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(wr_data[7]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(wr_data[8]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(wr_data[9]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(wr_valid),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(cmd_ready));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(init_done));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(phy_addr[0]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net105),
    .X(phy_addr[10]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net106),
    .X(phy_addr[11]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net107),
    .X(phy_addr[12]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net108),
    .X(phy_addr[13]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net109),
    .X(phy_addr[1]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net110),
    .X(phy_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net111),
    .X(phy_addr[3]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net112),
    .X(phy_addr[4]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net113),
    .X(phy_addr[5]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net114),
    .X(phy_addr[6]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net115),
    .X(phy_addr[7]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net116),
    .X(phy_addr[8]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net117),
    .X(phy_addr[9]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net118),
    .X(phy_bank[0]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net119),
    .X(phy_bank[1]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net120),
    .X(phy_bank[2]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net121),
    .X(phy_cas_n));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net122),
    .X(phy_cs_n));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net123),
    .X(phy_dm[0]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net124),
    .X(phy_dm[1]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net125),
    .X(phy_dm[2]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net126),
    .X(phy_dm[3]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net127),
    .X(phy_dm[4]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net128),
    .X(phy_dm[5]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net129),
    .X(phy_dm[6]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net130),
    .X(phy_dm[7]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net131),
    .X(phy_ras_n));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net132),
    .X(phy_reset_n));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net133),
    .X(phy_we_n));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net134),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net135),
    .X(rd_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net136),
    .X(rd_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net137),
    .X(rd_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net138),
    .X(rd_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net139),
    .X(rd_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net140),
    .X(rd_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net141),
    .X(rd_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net142),
    .X(rd_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net143),
    .X(rd_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net144),
    .X(rd_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net145),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net146),
    .X(rd_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net147),
    .X(rd_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net148),
    .X(rd_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net149),
    .X(rd_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net150),
    .X(rd_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net151),
    .X(rd_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net152),
    .X(rd_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net153),
    .X(rd_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net154),
    .X(rd_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net155),
    .X(rd_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net156),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net157),
    .X(rd_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net158),
    .X(rd_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net159),
    .X(rd_data[32]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net160),
    .X(rd_data[33]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net161),
    .X(rd_data[34]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net162),
    .X(rd_data[35]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net163),
    .X(rd_data[36]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net164),
    .X(rd_data[37]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net165),
    .X(rd_data[38]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net166),
    .X(rd_data[39]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net167),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net168),
    .X(rd_data[40]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net169),
    .X(rd_data[41]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net170),
    .X(rd_data[42]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net171),
    .X(rd_data[43]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net172),
    .X(rd_data[44]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net173),
    .X(rd_data[45]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net174),
    .X(rd_data[46]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net175),
    .X(rd_data[47]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net176),
    .X(rd_data[48]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net177),
    .X(rd_data[49]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net178),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net179),
    .X(rd_data[50]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net180),
    .X(rd_data[51]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net181),
    .X(rd_data[52]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net182),
    .X(rd_data[53]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net183),
    .X(rd_data[54]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net184),
    .X(rd_data[55]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net185),
    .X(rd_data[56]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net186),
    .X(rd_data[57]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net187),
    .X(rd_data[58]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net188),
    .X(rd_data[59]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net189),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net190),
    .X(rd_data[60]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net191),
    .X(rd_data[61]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net192),
    .X(rd_data[62]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net193),
    .X(rd_data[63]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net194),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net195),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net196),
    .X(rd_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net197),
    .X(rd_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net198),
    .X(rd_valid));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net199),
    .X(state[0]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net200),
    .X(state[1]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net201),
    .X(wr_ready));
 sky130_fd_sc_hd__conb_1 _1326__201 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _1327__202 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _1401__203 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _1402__204 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _1403__205 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _1404__206 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _1405__207 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _1406__208 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _1407__209 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _1408__210 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _1409__212 (.HI(net213));
 sky130_fd_sc_hd__conb_1 _1410__213 (.HI(net214));
 sky130_fd_sc_hd__conb_1 _1411__214 (.HI(net215));
 sky130_fd_sc_hd__conb_1 _1412__215 (.HI(net216));
 sky130_fd_sc_hd__conb_1 _1413__216 (.HI(net217));
 sky130_fd_sc_hd__conb_1 _1414__217 (.HI(net218));
 sky130_fd_sc_hd__conb_1 _1415__218 (.HI(net219));
 sky130_fd_sc_hd__conb_1 _1416__219 (.HI(net220));
 sky130_fd_sc_hd__conb_1 _1417__220 (.HI(net221));
 sky130_fd_sc_hd__conb_1 \cmd_reg_valid$_DFF_PN0__221  (.HI(net222));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_8 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net223));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_298 ();
endmodule
