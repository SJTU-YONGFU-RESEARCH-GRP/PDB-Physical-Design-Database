module leading_zero_counter (valid_input,
    data_in,
    zero_count);
 output valid_input;
 input [31:0] data_in;
 output [5:0] zero_count;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;

 gf180mcu_fd_sc_mcu9t5v0__or2_2 _061_ (.A1(net32),
    .A2(net31),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _062_ (.A1(net3),
    .A2(net2),
    .A3(_006_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _063_ (.A1(net5),
    .A2(net4),
    .A3(net7),
    .A4(net6),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _064_ (.A1(net30),
    .A2(net29),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _065_ (.A1(net26),
    .A2(net23),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _066_ (.A1(net12),
    .A2(net1),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _067_ (.A1(net28),
    .A2(net27),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _068_ (.A1(_009_),
    .A2(_010_),
    .A3(_011_),
    .A4(_012_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _069_ (.I(_013_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _070_ (.A1(_007_),
    .A2(_008_),
    .A3(_014_),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _071_ (.I(net9),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _072_ (.I(net8),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _073_ (.A1(net11),
    .A2(net10),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _074_ (.A1(net14),
    .A2(net13),
    .A3(net16),
    .A4(net15),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _075_ (.A1(_015_),
    .A2(_016_),
    .A3(_017_),
    .A4(_018_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _076_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net19),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _077_ (.A1(net22),
    .A2(net21),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _078_ (.A1(net25),
    .A2(net24),
    .A3(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _079_ (.A1(net38),
    .A2(_019_),
    .A3(_020_),
    .A4(_022_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _080_ (.A1(net38),
    .A2(_019_),
    .A3(_020_),
    .A4(_022_),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _081_ (.I(net19),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _082_ (.I(net22),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _083_ (.A1(_024_),
    .A2(net24),
    .B(net21),
    .C(net19),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _084_ (.A1(net20),
    .A2(_023_),
    .B(_025_),
    .C(net18),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _085_ (.A1(net13),
    .A2(net15),
    .A3(net17),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _086_ (.I(net13),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _087_ (.A1(net13),
    .A2(net15),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _088_ (.A1(net7),
    .A2(net9),
    .A3(net11),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _089_ (.A1(net14),
    .A2(_028_),
    .B1(net16),
    .B2(_029_),
    .C(_030_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _090_ (.A1(_026_),
    .A2(_027_),
    .B(_031_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _091_ (.I(net30),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _092_ (.A1(_033_),
    .A2(net31),
    .B(net29),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _093_ (.A1(net1),
    .A2(net23),
    .A3(net27),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _094_ (.A1(net28),
    .A2(_034_),
    .B(_035_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _095_ (.A1(_015_),
    .A2(net10),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _096_ (.A1(_016_),
    .A2(_037_),
    .B(net7),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _097_ (.A1(net2),
    .A2(net4),
    .A3(net6),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _098_ (.A1(_036_),
    .A2(_038_),
    .A3(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _099_ (.I(net4),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _100_ (.A1(net5),
    .A2(_041_),
    .B(net3),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _101_ (.A1(net2),
    .A2(_042_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _102_ (.A1(net28),
    .A2(net30),
    .A3(net32),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _103_ (.A1(_043_),
    .A2(_044_),
    .B(_036_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _104_ (.I(net23),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _105_ (.A1(net26),
    .A2(_046_),
    .B(net12),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _106_ (.A1(net1),
    .A2(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _107_ (.A1(_032_),
    .A2(_040_),
    .B(_045_),
    .C(_048_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _108_ (.A1(net20),
    .A2(net19),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _109_ (.A1(_049_),
    .A2(_021_),
    .B(net18),
    .C(net17),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _110_ (.A1(net14),
    .A2(net13),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _111_ (.A1(net16),
    .A2(net15),
    .A3(_050_),
    .B(_051_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _112_ (.A1(net5),
    .A2(net4),
    .A3(net9),
    .A4(net8),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _113_ (.A1(_017_),
    .A2(_052_),
    .B(_053_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _114_ (.A1(_009_),
    .A2(_010_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _115_ (.A1(net7),
    .A2(net6),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _116_ (.A1(net5),
    .A2(net4),
    .A3(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _117_ (.A1(net3),
    .A2(net2),
    .A3(_055_),
    .A4(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _118_ (.A1(_006_),
    .A2(_009_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _119_ (.A1(net28),
    .A2(net27),
    .A3(_059_),
    .B(_010_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _120_ (.A1(_054_),
    .A2(_058_),
    .B(_060_),
    .C(_011_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _121_ (.A1(_009_),
    .A2(_012_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _122_ (.A1(net9),
    .A2(net8),
    .A3(net11),
    .A4(net10),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _123_ (.A1(_018_),
    .A2(_020_),
    .B(_001_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _124_ (.A1(_008_),
    .A2(_002_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _125_ (.A1(_007_),
    .A2(_003_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _126_ (.A1(_000_),
    .A2(_004_),
    .B(_010_),
    .C(_011_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _127_ (.I(_019_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _128_ (.A1(_007_),
    .A2(_008_),
    .A3(_005_),
    .B(_013_),
    .ZN(net37));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_75 ();
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input1 (.I(data_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(data_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(data_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input4 (.I(data_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input5 (.I(data_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(data_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input7 (.I(data_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(data_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(data_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(data_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(data_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(data_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(data_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input14 (.I(data_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(data_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input16 (.I(data_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(data_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(data_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input19 (.I(data_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(data_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(data_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(data_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input23 (.I(data_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(data_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(data_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(data_in[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input27 (.I(data_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input28 (.I(data_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(data_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input30 (.I(data_in[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(data_in[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(data_in[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output33 (.I(net33),
    .Z(valid_input));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net34),
    .Z(zero_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net35),
    .Z(zero_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net36),
    .Z(zero_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net37),
    .Z(zero_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net38),
    .Z(zero_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net39),
    .Z(zero_count[5]));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_280 ();
endmodule
