module shadow_register (clk,
    main_load_en,
    rst_n,
    shadow_capture_en,
    shadow_load_en,
    use_shadow_out,
    main_data_in,
    main_data_out,
    shadow_data_in,
    shadow_data_out);
 input clk;
 input main_load_en;
 input rst_n;
 input shadow_capture_en;
 input shadow_load_en;
 input use_shadow_out;
 input [31:0] main_data_in;
 output [31:0] main_data_out;
 input [31:0] shadow_data_in;
 output [31:0] shadow_data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire \main_reg[0] ;
 wire \main_reg[10] ;
 wire \main_reg[11] ;
 wire \main_reg[12] ;
 wire \main_reg[13] ;
 wire \main_reg[14] ;
 wire \main_reg[15] ;
 wire \main_reg[16] ;
 wire \main_reg[17] ;
 wire \main_reg[18] ;
 wire \main_reg[19] ;
 wire \main_reg[1] ;
 wire \main_reg[20] ;
 wire \main_reg[21] ;
 wire \main_reg[22] ;
 wire \main_reg[23] ;
 wire \main_reg[24] ;
 wire \main_reg[25] ;
 wire \main_reg[26] ;
 wire \main_reg[27] ;
 wire \main_reg[28] ;
 wire \main_reg[29] ;
 wire \main_reg[2] ;
 wire \main_reg[30] ;
 wire \main_reg[31] ;
 wire \main_reg[3] ;
 wire \main_reg[4] ;
 wire \main_reg[5] ;
 wire \main_reg[6] ;
 wire \main_reg[7] ;
 wire \main_reg[8] ;
 wire \main_reg[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 CLKBUF_X3 _247_ (.A(rst_n),
    .Z(_064_));
 BUF_X2 _248_ (.A(_064_),
    .Z(_065_));
 BUF_X2 _249_ (.A(main_load_en),
    .Z(_066_));
 BUF_X4 _250_ (.A(_066_),
    .Z(_067_));
 MUX2_X1 _251_ (.A(\main_reg[0] ),
    .B(net1),
    .S(_067_),
    .Z(_068_));
 AND2_X1 _252_ (.A1(_065_),
    .A2(_068_),
    .ZN(_000_));
 MUX2_X1 _253_ (.A(\main_reg[10] ),
    .B(net2),
    .S(_067_),
    .Z(_069_));
 AND2_X1 _254_ (.A1(_065_),
    .A2(_069_),
    .ZN(_001_));
 MUX2_X1 _255_ (.A(\main_reg[11] ),
    .B(net3),
    .S(_067_),
    .Z(_070_));
 AND2_X1 _256_ (.A1(_065_),
    .A2(_070_),
    .ZN(_002_));
 MUX2_X1 _257_ (.A(\main_reg[12] ),
    .B(net4),
    .S(_067_),
    .Z(_071_));
 AND2_X1 _258_ (.A1(_065_),
    .A2(_071_),
    .ZN(_003_));
 MUX2_X1 _259_ (.A(\main_reg[13] ),
    .B(net5),
    .S(_067_),
    .Z(_072_));
 AND2_X1 _260_ (.A1(_065_),
    .A2(_072_),
    .ZN(_004_));
 MUX2_X1 _261_ (.A(\main_reg[14] ),
    .B(net6),
    .S(_067_),
    .Z(_073_));
 AND2_X1 _262_ (.A1(_065_),
    .A2(_073_),
    .ZN(_005_));
 MUX2_X1 _263_ (.A(\main_reg[15] ),
    .B(net7),
    .S(_067_),
    .Z(_074_));
 AND2_X1 _264_ (.A1(_065_),
    .A2(_074_),
    .ZN(_006_));
 MUX2_X1 _265_ (.A(\main_reg[16] ),
    .B(net8),
    .S(_067_),
    .Z(_075_));
 AND2_X1 _266_ (.A1(_065_),
    .A2(_075_),
    .ZN(_007_));
 MUX2_X1 _267_ (.A(\main_reg[17] ),
    .B(net9),
    .S(_067_),
    .Z(_076_));
 AND2_X1 _268_ (.A1(_065_),
    .A2(_076_),
    .ZN(_008_));
 MUX2_X1 _269_ (.A(\main_reg[18] ),
    .B(net10),
    .S(_067_),
    .Z(_077_));
 AND2_X1 _270_ (.A1(_065_),
    .A2(_077_),
    .ZN(_009_));
 BUF_X2 _271_ (.A(_064_),
    .Z(_078_));
 BUF_X4 _272_ (.A(_066_),
    .Z(_079_));
 MUX2_X1 _273_ (.A(\main_reg[19] ),
    .B(net11),
    .S(_079_),
    .Z(_080_));
 AND2_X1 _274_ (.A1(_078_),
    .A2(_080_),
    .ZN(_010_));
 MUX2_X1 _275_ (.A(\main_reg[1] ),
    .B(net12),
    .S(_079_),
    .Z(_081_));
 AND2_X1 _276_ (.A1(_078_),
    .A2(_081_),
    .ZN(_011_));
 MUX2_X1 _277_ (.A(\main_reg[20] ),
    .B(net13),
    .S(_079_),
    .Z(_082_));
 AND2_X1 _278_ (.A1(_078_),
    .A2(_082_),
    .ZN(_012_));
 MUX2_X1 _279_ (.A(\main_reg[21] ),
    .B(net14),
    .S(_079_),
    .Z(_083_));
 AND2_X1 _280_ (.A1(_078_),
    .A2(_083_),
    .ZN(_013_));
 MUX2_X1 _281_ (.A(\main_reg[22] ),
    .B(net15),
    .S(_079_),
    .Z(_084_));
 AND2_X1 _282_ (.A1(_078_),
    .A2(_084_),
    .ZN(_014_));
 MUX2_X1 _283_ (.A(\main_reg[23] ),
    .B(net16),
    .S(_079_),
    .Z(_085_));
 AND2_X1 _284_ (.A1(_078_),
    .A2(_085_),
    .ZN(_015_));
 MUX2_X1 _285_ (.A(\main_reg[24] ),
    .B(net17),
    .S(_079_),
    .Z(_086_));
 AND2_X1 _286_ (.A1(_078_),
    .A2(_086_),
    .ZN(_016_));
 MUX2_X1 _287_ (.A(\main_reg[25] ),
    .B(net18),
    .S(_079_),
    .Z(_087_));
 AND2_X1 _288_ (.A1(_078_),
    .A2(_087_),
    .ZN(_017_));
 MUX2_X1 _289_ (.A(\main_reg[26] ),
    .B(net19),
    .S(_079_),
    .Z(_088_));
 AND2_X1 _290_ (.A1(_078_),
    .A2(_088_),
    .ZN(_018_));
 MUX2_X1 _291_ (.A(\main_reg[27] ),
    .B(net20),
    .S(_079_),
    .Z(_089_));
 AND2_X1 _292_ (.A1(_078_),
    .A2(_089_),
    .ZN(_019_));
 BUF_X2 _293_ (.A(_064_),
    .Z(_090_));
 BUF_X4 _294_ (.A(_066_),
    .Z(_091_));
 MUX2_X1 _295_ (.A(\main_reg[28] ),
    .B(net21),
    .S(_091_),
    .Z(_092_));
 AND2_X1 _296_ (.A1(_090_),
    .A2(_092_),
    .ZN(_020_));
 MUX2_X1 _297_ (.A(\main_reg[29] ),
    .B(net22),
    .S(_091_),
    .Z(_093_));
 AND2_X1 _298_ (.A1(_090_),
    .A2(_093_),
    .ZN(_021_));
 MUX2_X1 _299_ (.A(\main_reg[2] ),
    .B(net23),
    .S(_091_),
    .Z(_094_));
 AND2_X1 _300_ (.A1(_090_),
    .A2(_094_),
    .ZN(_022_));
 MUX2_X1 _301_ (.A(\main_reg[30] ),
    .B(net24),
    .S(_091_),
    .Z(_095_));
 AND2_X1 _302_ (.A1(_090_),
    .A2(_095_),
    .ZN(_023_));
 MUX2_X1 _303_ (.A(\main_reg[31] ),
    .B(net25),
    .S(_091_),
    .Z(_096_));
 AND2_X1 _304_ (.A1(_090_),
    .A2(_096_),
    .ZN(_024_));
 MUX2_X1 _305_ (.A(\main_reg[3] ),
    .B(net26),
    .S(_091_),
    .Z(_097_));
 AND2_X1 _306_ (.A1(_090_),
    .A2(_097_),
    .ZN(_025_));
 MUX2_X1 _307_ (.A(\main_reg[4] ),
    .B(net27),
    .S(_091_),
    .Z(_098_));
 AND2_X1 _308_ (.A1(_090_),
    .A2(_098_),
    .ZN(_026_));
 MUX2_X1 _309_ (.A(\main_reg[5] ),
    .B(net28),
    .S(_091_),
    .Z(_099_));
 AND2_X1 _310_ (.A1(_090_),
    .A2(_099_),
    .ZN(_027_));
 MUX2_X1 _311_ (.A(\main_reg[6] ),
    .B(net29),
    .S(_091_),
    .Z(_100_));
 AND2_X1 _312_ (.A1(_090_),
    .A2(_100_),
    .ZN(_028_));
 MUX2_X1 _313_ (.A(\main_reg[7] ),
    .B(net30),
    .S(_091_),
    .Z(_101_));
 AND2_X1 _314_ (.A1(_090_),
    .A2(_101_),
    .ZN(_029_));
 BUF_X2 _315_ (.A(_064_),
    .Z(_102_));
 MUX2_X1 _316_ (.A(\main_reg[8] ),
    .B(net31),
    .S(_066_),
    .Z(_103_));
 AND2_X1 _317_ (.A1(_102_),
    .A2(_103_),
    .ZN(_030_));
 MUX2_X1 _318_ (.A(\main_reg[9] ),
    .B(net32),
    .S(_066_),
    .Z(_104_));
 AND2_X1 _319_ (.A1(_102_),
    .A2(_104_),
    .ZN(_031_));
 BUF_X8 _320_ (.A(shadow_load_en),
    .Z(_105_));
 BUF_X8 _321_ (.A(_105_),
    .Z(_106_));
 MUX2_X1 _322_ (.A(net97),
    .B(net33),
    .S(_106_),
    .Z(_107_));
 CLKBUF_X3 _323_ (.A(shadow_capture_en),
    .Z(_108_));
 BUF_X4 _324_ (.A(_108_),
    .Z(_109_));
 MUX2_X1 _325_ (.A(_107_),
    .B(\main_reg[0] ),
    .S(_109_),
    .Z(_110_));
 AND2_X1 _326_ (.A1(_102_),
    .A2(_110_),
    .ZN(_032_));
 MUX2_X1 _327_ (.A(net98),
    .B(net34),
    .S(_106_),
    .Z(_111_));
 MUX2_X1 _328_ (.A(_111_),
    .B(\main_reg[10] ),
    .S(_109_),
    .Z(_112_));
 AND2_X1 _329_ (.A1(_102_),
    .A2(_112_),
    .ZN(_033_));
 MUX2_X1 _330_ (.A(net99),
    .B(net35),
    .S(_106_),
    .Z(_113_));
 MUX2_X1 _331_ (.A(_113_),
    .B(\main_reg[11] ),
    .S(_109_),
    .Z(_114_));
 AND2_X1 _332_ (.A1(_102_),
    .A2(_114_),
    .ZN(_034_));
 MUX2_X1 _333_ (.A(net100),
    .B(net36),
    .S(_106_),
    .Z(_115_));
 MUX2_X1 _334_ (.A(_115_),
    .B(\main_reg[12] ),
    .S(_109_),
    .Z(_116_));
 AND2_X1 _335_ (.A1(_102_),
    .A2(_116_),
    .ZN(_035_));
 MUX2_X1 _336_ (.A(net101),
    .B(net37),
    .S(_106_),
    .Z(_117_));
 MUX2_X1 _337_ (.A(_117_),
    .B(\main_reg[13] ),
    .S(_109_),
    .Z(_118_));
 AND2_X1 _338_ (.A1(_102_),
    .A2(_118_),
    .ZN(_036_));
 MUX2_X1 _339_ (.A(net102),
    .B(net38),
    .S(_106_),
    .Z(_119_));
 MUX2_X1 _340_ (.A(_119_),
    .B(\main_reg[14] ),
    .S(_109_),
    .Z(_120_));
 AND2_X1 _341_ (.A1(_102_),
    .A2(_120_),
    .ZN(_037_));
 MUX2_X1 _342_ (.A(net103),
    .B(net39),
    .S(_106_),
    .Z(_121_));
 MUX2_X1 _343_ (.A(_121_),
    .B(\main_reg[15] ),
    .S(_109_),
    .Z(_122_));
 AND2_X1 _344_ (.A1(_102_),
    .A2(_122_),
    .ZN(_038_));
 MUX2_X1 _345_ (.A(net104),
    .B(net40),
    .S(_106_),
    .Z(_123_));
 MUX2_X1 _346_ (.A(_123_),
    .B(\main_reg[16] ),
    .S(_109_),
    .Z(_124_));
 AND2_X1 _347_ (.A1(_102_),
    .A2(_124_),
    .ZN(_039_));
 BUF_X2 _348_ (.A(_064_),
    .Z(_125_));
 MUX2_X1 _349_ (.A(net105),
    .B(net41),
    .S(_106_),
    .Z(_126_));
 MUX2_X1 _350_ (.A(_126_),
    .B(\main_reg[17] ),
    .S(_109_),
    .Z(_127_));
 AND2_X1 _351_ (.A1(_125_),
    .A2(_127_),
    .ZN(_040_));
 MUX2_X1 _352_ (.A(net106),
    .B(net42),
    .S(_106_),
    .Z(_128_));
 MUX2_X1 _353_ (.A(_128_),
    .B(\main_reg[18] ),
    .S(_109_),
    .Z(_129_));
 AND2_X1 _354_ (.A1(_125_),
    .A2(_129_),
    .ZN(_041_));
 BUF_X8 _355_ (.A(_105_),
    .Z(_130_));
 MUX2_X1 _356_ (.A(net107),
    .B(net43),
    .S(_130_),
    .Z(_131_));
 BUF_X4 _357_ (.A(_108_),
    .Z(_132_));
 MUX2_X1 _358_ (.A(_131_),
    .B(\main_reg[19] ),
    .S(_132_),
    .Z(_133_));
 AND2_X1 _359_ (.A1(_125_),
    .A2(_133_),
    .ZN(_042_));
 MUX2_X1 _360_ (.A(net108),
    .B(net44),
    .S(_130_),
    .Z(_134_));
 MUX2_X1 _361_ (.A(_134_),
    .B(\main_reg[1] ),
    .S(_132_),
    .Z(_135_));
 AND2_X1 _362_ (.A1(_125_),
    .A2(_135_),
    .ZN(_043_));
 MUX2_X1 _363_ (.A(net109),
    .B(net45),
    .S(_130_),
    .Z(_136_));
 MUX2_X1 _364_ (.A(_136_),
    .B(\main_reg[20] ),
    .S(_132_),
    .Z(_137_));
 AND2_X1 _365_ (.A1(_125_),
    .A2(_137_),
    .ZN(_044_));
 MUX2_X1 _366_ (.A(net110),
    .B(net46),
    .S(_130_),
    .Z(_138_));
 MUX2_X1 _367_ (.A(_138_),
    .B(\main_reg[21] ),
    .S(_132_),
    .Z(_139_));
 AND2_X1 _368_ (.A1(_125_),
    .A2(_139_),
    .ZN(_045_));
 MUX2_X1 _369_ (.A(net111),
    .B(net47),
    .S(_130_),
    .Z(_140_));
 MUX2_X1 _370_ (.A(_140_),
    .B(\main_reg[22] ),
    .S(_132_),
    .Z(_141_));
 AND2_X1 _371_ (.A1(_125_),
    .A2(_141_),
    .ZN(_046_));
 MUX2_X1 _372_ (.A(net112),
    .B(net48),
    .S(_130_),
    .Z(_142_));
 MUX2_X1 _373_ (.A(_142_),
    .B(\main_reg[23] ),
    .S(_132_),
    .Z(_143_));
 AND2_X1 _374_ (.A1(_125_),
    .A2(_143_),
    .ZN(_047_));
 MUX2_X1 _375_ (.A(net113),
    .B(net49),
    .S(_130_),
    .Z(_144_));
 MUX2_X1 _376_ (.A(_144_),
    .B(\main_reg[24] ),
    .S(_132_),
    .Z(_145_));
 AND2_X1 _377_ (.A1(_125_),
    .A2(_145_),
    .ZN(_048_));
 MUX2_X1 _378_ (.A(net114),
    .B(net50),
    .S(_130_),
    .Z(_146_));
 MUX2_X1 _379_ (.A(_146_),
    .B(\main_reg[25] ),
    .S(_132_),
    .Z(_147_));
 AND2_X1 _380_ (.A1(_125_),
    .A2(_147_),
    .ZN(_049_));
 BUF_X2 _381_ (.A(_064_),
    .Z(_148_));
 MUX2_X1 _382_ (.A(net115),
    .B(net51),
    .S(_130_),
    .Z(_149_));
 MUX2_X1 _383_ (.A(_149_),
    .B(\main_reg[26] ),
    .S(_132_),
    .Z(_150_));
 AND2_X1 _384_ (.A1(_148_),
    .A2(_150_),
    .ZN(_050_));
 MUX2_X1 _385_ (.A(net116),
    .B(net52),
    .S(_130_),
    .Z(_151_));
 MUX2_X1 _386_ (.A(_151_),
    .B(\main_reg[27] ),
    .S(_132_),
    .Z(_152_));
 AND2_X1 _387_ (.A1(_148_),
    .A2(_152_),
    .ZN(_051_));
 BUF_X8 _388_ (.A(_105_),
    .Z(_153_));
 MUX2_X1 _389_ (.A(net117),
    .B(net53),
    .S(_153_),
    .Z(_154_));
 BUF_X4 _390_ (.A(_108_),
    .Z(_155_));
 MUX2_X1 _391_ (.A(_154_),
    .B(\main_reg[28] ),
    .S(_155_),
    .Z(_156_));
 AND2_X1 _392_ (.A1(_148_),
    .A2(_156_),
    .ZN(_052_));
 MUX2_X1 _393_ (.A(net118),
    .B(net54),
    .S(_153_),
    .Z(_157_));
 MUX2_X1 _394_ (.A(_157_),
    .B(\main_reg[29] ),
    .S(_155_),
    .Z(_158_));
 AND2_X1 _395_ (.A1(_148_),
    .A2(_158_),
    .ZN(_053_));
 MUX2_X1 _396_ (.A(net119),
    .B(net55),
    .S(_153_),
    .Z(_159_));
 MUX2_X1 _397_ (.A(_159_),
    .B(\main_reg[2] ),
    .S(_155_),
    .Z(_160_));
 AND2_X1 _398_ (.A1(_148_),
    .A2(_160_),
    .ZN(_054_));
 MUX2_X1 _399_ (.A(net120),
    .B(net56),
    .S(_153_),
    .Z(_161_));
 MUX2_X1 _400_ (.A(_161_),
    .B(\main_reg[30] ),
    .S(_155_),
    .Z(_162_));
 AND2_X1 _401_ (.A1(_148_),
    .A2(_162_),
    .ZN(_055_));
 MUX2_X1 _402_ (.A(net121),
    .B(net57),
    .S(_153_),
    .Z(_163_));
 MUX2_X1 _403_ (.A(_163_),
    .B(\main_reg[31] ),
    .S(_155_),
    .Z(_164_));
 AND2_X1 _404_ (.A1(_148_),
    .A2(_164_),
    .ZN(_056_));
 MUX2_X1 _405_ (.A(net122),
    .B(net58),
    .S(_153_),
    .Z(_165_));
 MUX2_X1 _406_ (.A(_165_),
    .B(\main_reg[3] ),
    .S(_155_),
    .Z(_166_));
 AND2_X1 _407_ (.A1(_148_),
    .A2(_166_),
    .ZN(_057_));
 MUX2_X1 _408_ (.A(net123),
    .B(net59),
    .S(_153_),
    .Z(_167_));
 MUX2_X1 _409_ (.A(_167_),
    .B(\main_reg[4] ),
    .S(_155_),
    .Z(_168_));
 AND2_X1 _410_ (.A1(_148_),
    .A2(_168_),
    .ZN(_058_));
 MUX2_X1 _411_ (.A(net124),
    .B(net60),
    .S(_153_),
    .Z(_169_));
 MUX2_X1 _412_ (.A(_169_),
    .B(\main_reg[5] ),
    .S(_155_),
    .Z(_170_));
 AND2_X1 _413_ (.A1(_148_),
    .A2(_170_),
    .ZN(_059_));
 MUX2_X1 _414_ (.A(net125),
    .B(net61),
    .S(_153_),
    .Z(_171_));
 MUX2_X1 _415_ (.A(_171_),
    .B(\main_reg[6] ),
    .S(_155_),
    .Z(_172_));
 AND2_X1 _416_ (.A1(_064_),
    .A2(_172_),
    .ZN(_060_));
 MUX2_X1 _417_ (.A(net126),
    .B(net62),
    .S(_153_),
    .Z(_173_));
 MUX2_X1 _418_ (.A(_173_),
    .B(\main_reg[7] ),
    .S(_155_),
    .Z(_174_));
 AND2_X1 _419_ (.A1(_064_),
    .A2(_174_),
    .ZN(_061_));
 MUX2_X1 _420_ (.A(net127),
    .B(net63),
    .S(_105_),
    .Z(_175_));
 MUX2_X1 _421_ (.A(_175_),
    .B(\main_reg[8] ),
    .S(_108_),
    .Z(_176_));
 AND2_X1 _422_ (.A1(_064_),
    .A2(_176_),
    .ZN(_062_));
 MUX2_X1 _423_ (.A(net128),
    .B(net64),
    .S(_105_),
    .Z(_177_));
 MUX2_X1 _424_ (.A(_177_),
    .B(\main_reg[9] ),
    .S(_108_),
    .Z(_178_));
 AND2_X1 _425_ (.A1(_064_),
    .A2(_178_),
    .ZN(_063_));
 CLKBUF_X3 _426_ (.A(use_shadow_out),
    .Z(_179_));
 BUF_X4 _427_ (.A(_179_),
    .Z(_180_));
 MUX2_X1 _428_ (.A(\main_reg[0] ),
    .B(net97),
    .S(_180_),
    .Z(net65));
 MUX2_X1 _429_ (.A(\main_reg[10] ),
    .B(net98),
    .S(_180_),
    .Z(net66));
 MUX2_X1 _430_ (.A(\main_reg[11] ),
    .B(net99),
    .S(_180_),
    .Z(net67));
 MUX2_X1 _431_ (.A(\main_reg[12] ),
    .B(net100),
    .S(_180_),
    .Z(net68));
 MUX2_X1 _432_ (.A(\main_reg[13] ),
    .B(net101),
    .S(_180_),
    .Z(net69));
 MUX2_X1 _433_ (.A(\main_reg[14] ),
    .B(net102),
    .S(_180_),
    .Z(net70));
 MUX2_X1 _434_ (.A(\main_reg[15] ),
    .B(net103),
    .S(_180_),
    .Z(net71));
 MUX2_X1 _435_ (.A(\main_reg[16] ),
    .B(net104),
    .S(_180_),
    .Z(net72));
 MUX2_X1 _436_ (.A(\main_reg[17] ),
    .B(net105),
    .S(_180_),
    .Z(net73));
 MUX2_X1 _437_ (.A(\main_reg[18] ),
    .B(net106),
    .S(_180_),
    .Z(net74));
 BUF_X4 _438_ (.A(_179_),
    .Z(_181_));
 MUX2_X1 _439_ (.A(\main_reg[19] ),
    .B(net107),
    .S(_181_),
    .Z(net75));
 MUX2_X1 _440_ (.A(\main_reg[1] ),
    .B(net108),
    .S(_181_),
    .Z(net76));
 MUX2_X1 _441_ (.A(\main_reg[20] ),
    .B(net109),
    .S(_181_),
    .Z(net77));
 MUX2_X1 _442_ (.A(\main_reg[21] ),
    .B(net110),
    .S(_181_),
    .Z(net78));
 MUX2_X1 _443_ (.A(\main_reg[22] ),
    .B(net111),
    .S(_181_),
    .Z(net79));
 MUX2_X1 _444_ (.A(\main_reg[23] ),
    .B(net112),
    .S(_181_),
    .Z(net80));
 MUX2_X1 _445_ (.A(\main_reg[24] ),
    .B(net113),
    .S(_181_),
    .Z(net81));
 MUX2_X1 _446_ (.A(\main_reg[25] ),
    .B(net114),
    .S(_181_),
    .Z(net82));
 MUX2_X1 _447_ (.A(\main_reg[26] ),
    .B(net115),
    .S(_181_),
    .Z(net83));
 MUX2_X1 _448_ (.A(\main_reg[27] ),
    .B(net116),
    .S(_181_),
    .Z(net84));
 BUF_X4 _449_ (.A(_179_),
    .Z(_182_));
 MUX2_X1 _450_ (.A(\main_reg[28] ),
    .B(net117),
    .S(_182_),
    .Z(net85));
 MUX2_X1 _451_ (.A(\main_reg[29] ),
    .B(net118),
    .S(_182_),
    .Z(net86));
 MUX2_X1 _452_ (.A(\main_reg[2] ),
    .B(net119),
    .S(_182_),
    .Z(net87));
 MUX2_X1 _453_ (.A(\main_reg[30] ),
    .B(net120),
    .S(_182_),
    .Z(net88));
 MUX2_X1 _454_ (.A(\main_reg[31] ),
    .B(net121),
    .S(_182_),
    .Z(net89));
 MUX2_X1 _455_ (.A(\main_reg[3] ),
    .B(net122),
    .S(_182_),
    .Z(net90));
 MUX2_X1 _456_ (.A(\main_reg[4] ),
    .B(net123),
    .S(_182_),
    .Z(net91));
 MUX2_X1 _457_ (.A(\main_reg[5] ),
    .B(net124),
    .S(_182_),
    .Z(net92));
 MUX2_X1 _458_ (.A(\main_reg[6] ),
    .B(net125),
    .S(_182_),
    .Z(net93));
 MUX2_X1 _459_ (.A(\main_reg[7] ),
    .B(net126),
    .S(_182_),
    .Z(net94));
 MUX2_X1 _460_ (.A(\main_reg[8] ),
    .B(net127),
    .S(_179_),
    .Z(net95));
 MUX2_X1 _461_ (.A(\main_reg[9] ),
    .B(net128),
    .S(_179_),
    .Z(net96));
 DFF_X1 \main_reg[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\main_reg[0] ),
    .QN(_246_));
 DFF_X1 \main_reg[10]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\main_reg[10] ),
    .QN(_245_));
 DFF_X1 \main_reg[11]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\main_reg[11] ),
    .QN(_244_));
 DFF_X1 \main_reg[12]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\main_reg[12] ),
    .QN(_243_));
 DFF_X1 \main_reg[13]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\main_reg[13] ),
    .QN(_242_));
 DFF_X1 \main_reg[14]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\main_reg[14] ),
    .QN(_241_));
 DFF_X1 \main_reg[15]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\main_reg[15] ),
    .QN(_240_));
 DFF_X1 \main_reg[16]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\main_reg[16] ),
    .QN(_239_));
 DFF_X1 \main_reg[17]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\main_reg[17] ),
    .QN(_238_));
 DFF_X1 \main_reg[18]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\main_reg[18] ),
    .QN(_237_));
 DFF_X1 \main_reg[19]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\main_reg[19] ),
    .QN(_236_));
 DFF_X1 \main_reg[1]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\main_reg[1] ),
    .QN(_235_));
 DFF_X1 \main_reg[20]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\main_reg[20] ),
    .QN(_234_));
 DFF_X1 \main_reg[21]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\main_reg[21] ),
    .QN(_233_));
 DFF_X1 \main_reg[22]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\main_reg[22] ),
    .QN(_232_));
 DFF_X1 \main_reg[23]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\main_reg[23] ),
    .QN(_231_));
 DFF_X1 \main_reg[24]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\main_reg[24] ),
    .QN(_230_));
 DFF_X1 \main_reg[25]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\main_reg[25] ),
    .QN(_229_));
 DFF_X1 \main_reg[26]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\main_reg[26] ),
    .QN(_228_));
 DFF_X1 \main_reg[27]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\main_reg[27] ),
    .QN(_227_));
 DFF_X1 \main_reg[28]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\main_reg[28] ),
    .QN(_226_));
 DFF_X1 \main_reg[29]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\main_reg[29] ),
    .QN(_225_));
 DFF_X1 \main_reg[2]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\main_reg[2] ),
    .QN(_224_));
 DFF_X1 \main_reg[30]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\main_reg[30] ),
    .QN(_223_));
 DFF_X1 \main_reg[31]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\main_reg[31] ),
    .QN(_222_));
 DFF_X1 \main_reg[3]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\main_reg[3] ),
    .QN(_221_));
 DFF_X1 \main_reg[4]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\main_reg[4] ),
    .QN(_220_));
 DFF_X1 \main_reg[5]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\main_reg[5] ),
    .QN(_219_));
 DFF_X1 \main_reg[6]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\main_reg[6] ),
    .QN(_218_));
 DFF_X1 \main_reg[7]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\main_reg[7] ),
    .QN(_217_));
 DFF_X1 \main_reg[8]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\main_reg[8] ),
    .QN(_216_));
 DFF_X1 \main_reg[9]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\main_reg[9] ),
    .QN(_215_));
 DFF_X1 \shadow_reg[0]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net97),
    .QN(_214_));
 DFF_X1 \shadow_reg[10]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net98),
    .QN(_213_));
 DFF_X1 \shadow_reg[11]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net99),
    .QN(_212_));
 DFF_X1 \shadow_reg[12]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net100),
    .QN(_211_));
 DFF_X1 \shadow_reg[13]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net101),
    .QN(_210_));
 DFF_X1 \shadow_reg[14]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net102),
    .QN(_209_));
 DFF_X1 \shadow_reg[15]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net103),
    .QN(_208_));
 DFF_X1 \shadow_reg[16]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net104),
    .QN(_207_));
 DFF_X1 \shadow_reg[17]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net105),
    .QN(_206_));
 DFF_X1 \shadow_reg[18]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net106),
    .QN(_205_));
 DFF_X1 \shadow_reg[19]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net107),
    .QN(_204_));
 DFF_X1 \shadow_reg[1]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net108),
    .QN(_203_));
 DFF_X1 \shadow_reg[20]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net109),
    .QN(_202_));
 DFF_X1 \shadow_reg[21]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net110),
    .QN(_201_));
 DFF_X1 \shadow_reg[22]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net111),
    .QN(_200_));
 DFF_X1 \shadow_reg[23]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net112),
    .QN(_199_));
 DFF_X1 \shadow_reg[24]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net113),
    .QN(_198_));
 DFF_X1 \shadow_reg[25]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net114),
    .QN(_197_));
 DFF_X1 \shadow_reg[26]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net115),
    .QN(_196_));
 DFF_X1 \shadow_reg[27]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net116),
    .QN(_195_));
 DFF_X1 \shadow_reg[28]$_SDFFE_PN0P_  (.D(_052_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net117),
    .QN(_194_));
 DFF_X1 \shadow_reg[29]$_SDFFE_PN0P_  (.D(_053_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net118),
    .QN(_193_));
 DFF_X1 \shadow_reg[2]$_SDFFE_PN0P_  (.D(_054_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net119),
    .QN(_192_));
 DFF_X1 \shadow_reg[30]$_SDFFE_PN0P_  (.D(_055_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net120),
    .QN(_191_));
 DFF_X1 \shadow_reg[31]$_SDFFE_PN0P_  (.D(_056_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net121),
    .QN(_190_));
 DFF_X1 \shadow_reg[3]$_SDFFE_PN0P_  (.D(_057_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net122),
    .QN(_189_));
 DFF_X1 \shadow_reg[4]$_SDFFE_PN0P_  (.D(_058_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net123),
    .QN(_188_));
 DFF_X1 \shadow_reg[5]$_SDFFE_PN0P_  (.D(_059_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net124),
    .QN(_187_));
 DFF_X1 \shadow_reg[6]$_SDFFE_PN0P_  (.D(_060_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net125),
    .QN(_186_));
 DFF_X1 \shadow_reg[7]$_SDFFE_PN0P_  (.D(_061_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net126),
    .QN(_185_));
 DFF_X1 \shadow_reg[8]$_SDFFE_PN0P_  (.D(_062_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net127),
    .QN(_184_));
 DFF_X1 \shadow_reg[9]$_SDFFE_PN0P_  (.D(_063_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net128),
    .QN(_183_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_93 ();
 BUF_X1 input1 (.A(main_data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(main_data_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(main_data_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(main_data_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(main_data_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(main_data_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(main_data_in[15]),
    .Z(net7));
 BUF_X1 input8 (.A(main_data_in[16]),
    .Z(net8));
 BUF_X1 input9 (.A(main_data_in[17]),
    .Z(net9));
 BUF_X1 input10 (.A(main_data_in[18]),
    .Z(net10));
 BUF_X1 input11 (.A(main_data_in[19]),
    .Z(net11));
 BUF_X1 input12 (.A(main_data_in[1]),
    .Z(net12));
 BUF_X1 input13 (.A(main_data_in[20]),
    .Z(net13));
 BUF_X1 input14 (.A(main_data_in[21]),
    .Z(net14));
 BUF_X1 input15 (.A(main_data_in[22]),
    .Z(net15));
 BUF_X1 input16 (.A(main_data_in[23]),
    .Z(net16));
 BUF_X1 input17 (.A(main_data_in[24]),
    .Z(net17));
 BUF_X1 input18 (.A(main_data_in[25]),
    .Z(net18));
 BUF_X1 input19 (.A(main_data_in[26]),
    .Z(net19));
 BUF_X1 input20 (.A(main_data_in[27]),
    .Z(net20));
 BUF_X1 input21 (.A(main_data_in[28]),
    .Z(net21));
 BUF_X1 input22 (.A(main_data_in[29]),
    .Z(net22));
 BUF_X1 input23 (.A(main_data_in[2]),
    .Z(net23));
 BUF_X1 input24 (.A(main_data_in[30]),
    .Z(net24));
 BUF_X1 input25 (.A(main_data_in[31]),
    .Z(net25));
 BUF_X1 input26 (.A(main_data_in[3]),
    .Z(net26));
 BUF_X1 input27 (.A(main_data_in[4]),
    .Z(net27));
 BUF_X1 input28 (.A(main_data_in[5]),
    .Z(net28));
 BUF_X1 input29 (.A(main_data_in[6]),
    .Z(net29));
 BUF_X1 input30 (.A(main_data_in[7]),
    .Z(net30));
 BUF_X1 input31 (.A(main_data_in[8]),
    .Z(net31));
 BUF_X1 input32 (.A(main_data_in[9]),
    .Z(net32));
 BUF_X1 input33 (.A(shadow_data_in[0]),
    .Z(net33));
 BUF_X1 input34 (.A(shadow_data_in[10]),
    .Z(net34));
 BUF_X1 input35 (.A(shadow_data_in[11]),
    .Z(net35));
 BUF_X1 input36 (.A(shadow_data_in[12]),
    .Z(net36));
 BUF_X1 input37 (.A(shadow_data_in[13]),
    .Z(net37));
 BUF_X1 input38 (.A(shadow_data_in[14]),
    .Z(net38));
 BUF_X1 input39 (.A(shadow_data_in[15]),
    .Z(net39));
 BUF_X1 input40 (.A(shadow_data_in[16]),
    .Z(net40));
 BUF_X1 input41 (.A(shadow_data_in[17]),
    .Z(net41));
 BUF_X1 input42 (.A(shadow_data_in[18]),
    .Z(net42));
 BUF_X1 input43 (.A(shadow_data_in[19]),
    .Z(net43));
 BUF_X1 input44 (.A(shadow_data_in[1]),
    .Z(net44));
 BUF_X1 input45 (.A(shadow_data_in[20]),
    .Z(net45));
 BUF_X1 input46 (.A(shadow_data_in[21]),
    .Z(net46));
 BUF_X1 input47 (.A(shadow_data_in[22]),
    .Z(net47));
 BUF_X1 input48 (.A(shadow_data_in[23]),
    .Z(net48));
 BUF_X1 input49 (.A(shadow_data_in[24]),
    .Z(net49));
 BUF_X1 input50 (.A(shadow_data_in[25]),
    .Z(net50));
 BUF_X1 input51 (.A(shadow_data_in[26]),
    .Z(net51));
 BUF_X1 input52 (.A(shadow_data_in[27]),
    .Z(net52));
 BUF_X1 input53 (.A(shadow_data_in[28]),
    .Z(net53));
 BUF_X1 input54 (.A(shadow_data_in[29]),
    .Z(net54));
 BUF_X1 input55 (.A(shadow_data_in[2]),
    .Z(net55));
 BUF_X1 input56 (.A(shadow_data_in[30]),
    .Z(net56));
 BUF_X1 input57 (.A(shadow_data_in[31]),
    .Z(net57));
 BUF_X1 input58 (.A(shadow_data_in[3]),
    .Z(net58));
 BUF_X1 input59 (.A(shadow_data_in[4]),
    .Z(net59));
 BUF_X1 input60 (.A(shadow_data_in[5]),
    .Z(net60));
 BUF_X1 input61 (.A(shadow_data_in[6]),
    .Z(net61));
 BUF_X1 input62 (.A(shadow_data_in[7]),
    .Z(net62));
 BUF_X1 input63 (.A(shadow_data_in[8]),
    .Z(net63));
 BUF_X1 input64 (.A(shadow_data_in[9]),
    .Z(net64));
 BUF_X1 output65 (.A(net65),
    .Z(main_data_out[0]));
 BUF_X1 output66 (.A(net66),
    .Z(main_data_out[10]));
 BUF_X1 output67 (.A(net67),
    .Z(main_data_out[11]));
 BUF_X1 output68 (.A(net68),
    .Z(main_data_out[12]));
 BUF_X1 output69 (.A(net69),
    .Z(main_data_out[13]));
 BUF_X1 output70 (.A(net70),
    .Z(main_data_out[14]));
 BUF_X1 output71 (.A(net71),
    .Z(main_data_out[15]));
 BUF_X1 output72 (.A(net72),
    .Z(main_data_out[16]));
 BUF_X1 output73 (.A(net73),
    .Z(main_data_out[17]));
 BUF_X1 output74 (.A(net74),
    .Z(main_data_out[18]));
 BUF_X1 output75 (.A(net75),
    .Z(main_data_out[19]));
 BUF_X1 output76 (.A(net76),
    .Z(main_data_out[1]));
 BUF_X1 output77 (.A(net77),
    .Z(main_data_out[20]));
 BUF_X1 output78 (.A(net78),
    .Z(main_data_out[21]));
 BUF_X1 output79 (.A(net79),
    .Z(main_data_out[22]));
 BUF_X1 output80 (.A(net80),
    .Z(main_data_out[23]));
 BUF_X1 output81 (.A(net81),
    .Z(main_data_out[24]));
 BUF_X1 output82 (.A(net82),
    .Z(main_data_out[25]));
 BUF_X1 output83 (.A(net83),
    .Z(main_data_out[26]));
 BUF_X1 output84 (.A(net84),
    .Z(main_data_out[27]));
 BUF_X1 output85 (.A(net85),
    .Z(main_data_out[28]));
 BUF_X1 output86 (.A(net86),
    .Z(main_data_out[29]));
 BUF_X1 output87 (.A(net87),
    .Z(main_data_out[2]));
 BUF_X1 output88 (.A(net88),
    .Z(main_data_out[30]));
 BUF_X1 output89 (.A(net89),
    .Z(main_data_out[31]));
 BUF_X1 output90 (.A(net90),
    .Z(main_data_out[3]));
 BUF_X1 output91 (.A(net91),
    .Z(main_data_out[4]));
 BUF_X1 output92 (.A(net92),
    .Z(main_data_out[5]));
 BUF_X1 output93 (.A(net93),
    .Z(main_data_out[6]));
 BUF_X1 output94 (.A(net94),
    .Z(main_data_out[7]));
 BUF_X1 output95 (.A(net95),
    .Z(main_data_out[8]));
 BUF_X1 output96 (.A(net96),
    .Z(main_data_out[9]));
 BUF_X1 output97 (.A(net97),
    .Z(shadow_data_out[0]));
 BUF_X1 output98 (.A(net98),
    .Z(shadow_data_out[10]));
 BUF_X1 output99 (.A(net99),
    .Z(shadow_data_out[11]));
 BUF_X1 output100 (.A(net100),
    .Z(shadow_data_out[12]));
 BUF_X1 output101 (.A(net101),
    .Z(shadow_data_out[13]));
 BUF_X1 output102 (.A(net102),
    .Z(shadow_data_out[14]));
 BUF_X1 output103 (.A(net103),
    .Z(shadow_data_out[15]));
 BUF_X1 output104 (.A(net104),
    .Z(shadow_data_out[16]));
 BUF_X1 output105 (.A(net105),
    .Z(shadow_data_out[17]));
 BUF_X1 output106 (.A(net106),
    .Z(shadow_data_out[18]));
 BUF_X1 output107 (.A(net107),
    .Z(shadow_data_out[19]));
 BUF_X1 output108 (.A(net108),
    .Z(shadow_data_out[1]));
 BUF_X1 output109 (.A(net109),
    .Z(shadow_data_out[20]));
 BUF_X1 output110 (.A(net110),
    .Z(shadow_data_out[21]));
 BUF_X1 output111 (.A(net111),
    .Z(shadow_data_out[22]));
 BUF_X1 output112 (.A(net112),
    .Z(shadow_data_out[23]));
 BUF_X1 output113 (.A(net113),
    .Z(shadow_data_out[24]));
 BUF_X1 output114 (.A(net114),
    .Z(shadow_data_out[25]));
 BUF_X1 output115 (.A(net115),
    .Z(shadow_data_out[26]));
 BUF_X1 output116 (.A(net116),
    .Z(shadow_data_out[27]));
 BUF_X1 output117 (.A(net117),
    .Z(shadow_data_out[28]));
 BUF_X1 output118 (.A(net118),
    .Z(shadow_data_out[29]));
 BUF_X1 output119 (.A(net119),
    .Z(shadow_data_out[2]));
 BUF_X1 output120 (.A(net120),
    .Z(shadow_data_out[30]));
 BUF_X1 output121 (.A(net121),
    .Z(shadow_data_out[31]));
 BUF_X1 output122 (.A(net122),
    .Z(shadow_data_out[3]));
 BUF_X1 output123 (.A(net123),
    .Z(shadow_data_out[4]));
 BUF_X1 output124 (.A(net124),
    .Z(shadow_data_out[5]));
 BUF_X1 output125 (.A(net125),
    .Z(shadow_data_out[6]));
 BUF_X1 output126 (.A(net126),
    .Z(shadow_data_out[7]));
 BUF_X1 output127 (.A(net127),
    .Z(shadow_data_out[8]));
 BUF_X1 output128 (.A(net128),
    .Z(shadow_data_out[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X2 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X1 clkload2 (.A(clknet_3_3__leaf_clk));
 INV_X1 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_6__leaf_clk));
 CLKBUF_X1 clkload5 (.A(clknet_3_7__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_129 ();
 FILLCELL_X2 FILLER_0_133 ();
 FILLCELL_X1 FILLER_0_135 ();
 FILLCELL_X2 FILLER_0_151 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X2 FILLER_0_166 ();
 FILLCELL_X8 FILLER_0_171 ();
 FILLCELL_X4 FILLER_0_179 ();
 FILLCELL_X2 FILLER_0_183 ();
 FILLCELL_X1 FILLER_0_185 ();
 FILLCELL_X2 FILLER_0_195 ();
 FILLCELL_X8 FILLER_0_206 ();
 FILLCELL_X8 FILLER_0_217 ();
 FILLCELL_X4 FILLER_0_225 ();
 FILLCELL_X1 FILLER_0_229 ();
 FILLCELL_X4 FILLER_0_233 ();
 FILLCELL_X2 FILLER_0_237 ();
 FILLCELL_X2 FILLER_0_251 ();
 FILLCELL_X16 FILLER_0_256 ();
 FILLCELL_X2 FILLER_0_272 ();
 FILLCELL_X2 FILLER_0_277 ();
 FILLCELL_X1 FILLER_0_279 ();
 FILLCELL_X2 FILLER_0_286 ();
 FILLCELL_X1 FILLER_0_288 ();
 FILLCELL_X32 FILLER_0_292 ();
 FILLCELL_X16 FILLER_0_324 ();
 FILLCELL_X4 FILLER_0_340 ();
 FILLCELL_X2 FILLER_0_344 ();
 FILLCELL_X1 FILLER_0_346 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_97 ();
 FILLCELL_X8 FILLER_1_113 ();
 FILLCELL_X2 FILLER_1_121 ();
 FILLCELL_X1 FILLER_1_130 ();
 FILLCELL_X2 FILLER_1_138 ();
 FILLCELL_X4 FILLER_1_147 ();
 FILLCELL_X2 FILLER_1_151 ();
 FILLCELL_X1 FILLER_1_153 ();
 FILLCELL_X2 FILLER_1_164 ();
 FILLCELL_X2 FILLER_1_171 ();
 FILLCELL_X1 FILLER_1_173 ();
 FILLCELL_X1 FILLER_1_179 ();
 FILLCELL_X2 FILLER_1_193 ();
 FILLCELL_X1 FILLER_1_195 ();
 FILLCELL_X16 FILLER_1_206 ();
 FILLCELL_X8 FILLER_1_222 ();
 FILLCELL_X4 FILLER_1_230 ();
 FILLCELL_X2 FILLER_1_234 ();
 FILLCELL_X1 FILLER_1_236 ();
 FILLCELL_X8 FILLER_1_268 ();
 FILLCELL_X2 FILLER_1_276 ();
 FILLCELL_X32 FILLER_1_299 ();
 FILLCELL_X16 FILLER_1_331 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_97 ();
 FILLCELL_X2 FILLER_2_105 ();
 FILLCELL_X1 FILLER_2_107 ();
 FILLCELL_X8 FILLER_2_129 ();
 FILLCELL_X1 FILLER_2_137 ();
 FILLCELL_X2 FILLER_2_145 ();
 FILLCELL_X16 FILLER_2_168 ();
 FILLCELL_X4 FILLER_2_184 ();
 FILLCELL_X4 FILLER_2_220 ();
 FILLCELL_X2 FILLER_2_224 ();
 FILLCELL_X16 FILLER_2_233 ();
 FILLCELL_X8 FILLER_2_249 ();
 FILLCELL_X8 FILLER_2_261 ();
 FILLCELL_X4 FILLER_2_269 ();
 FILLCELL_X1 FILLER_2_273 ();
 FILLCELL_X32 FILLER_2_302 ();
 FILLCELL_X8 FILLER_2_334 ();
 FILLCELL_X4 FILLER_2_342 ();
 FILLCELL_X1 FILLER_2_346 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X16 FILLER_3_97 ();
 FILLCELL_X8 FILLER_3_113 ();
 FILLCELL_X1 FILLER_3_126 ();
 FILLCELL_X1 FILLER_3_152 ();
 FILLCELL_X16 FILLER_3_170 ();
 FILLCELL_X4 FILLER_3_186 ();
 FILLCELL_X2 FILLER_3_190 ();
 FILLCELL_X4 FILLER_3_209 ();
 FILLCELL_X2 FILLER_3_213 ();
 FILLCELL_X1 FILLER_3_215 ();
 FILLCELL_X8 FILLER_3_220 ();
 FILLCELL_X4 FILLER_3_228 ();
 FILLCELL_X8 FILLER_3_260 ();
 FILLCELL_X4 FILLER_3_268 ();
 FILLCELL_X1 FILLER_3_272 ();
 FILLCELL_X32 FILLER_3_294 ();
 FILLCELL_X16 FILLER_3_326 ();
 FILLCELL_X4 FILLER_3_342 ();
 FILLCELL_X1 FILLER_3_346 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X8 FILLER_4_193 ();
 FILLCELL_X4 FILLER_4_201 ();
 FILLCELL_X2 FILLER_4_205 ();
 FILLCELL_X32 FILLER_4_224 ();
 FILLCELL_X32 FILLER_4_256 ();
 FILLCELL_X32 FILLER_4_288 ();
 FILLCELL_X16 FILLER_4_320 ();
 FILLCELL_X8 FILLER_4_336 ();
 FILLCELL_X2 FILLER_4_344 ();
 FILLCELL_X1 FILLER_4_346 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X8 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_144 ();
 FILLCELL_X32 FILLER_5_176 ();
 FILLCELL_X32 FILLER_5_208 ();
 FILLCELL_X32 FILLER_5_240 ();
 FILLCELL_X4 FILLER_5_272 ();
 FILLCELL_X1 FILLER_5_276 ();
 FILLCELL_X32 FILLER_5_284 ();
 FILLCELL_X16 FILLER_5_316 ();
 FILLCELL_X8 FILLER_5_332 ();
 FILLCELL_X4 FILLER_5_340 ();
 FILLCELL_X2 FILLER_5_344 ();
 FILLCELL_X1 FILLER_5_346 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X8 FILLER_6_129 ();
 FILLCELL_X4 FILLER_6_137 ();
 FILLCELL_X8 FILLER_6_145 ();
 FILLCELL_X1 FILLER_6_153 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_177 ();
 FILLCELL_X2 FILLER_6_181 ();
 FILLCELL_X32 FILLER_6_221 ();
 FILLCELL_X16 FILLER_6_253 ();
 FILLCELL_X8 FILLER_6_269 ();
 FILLCELL_X4 FILLER_6_277 ();
 FILLCELL_X1 FILLER_6_281 ();
 FILLCELL_X32 FILLER_6_286 ();
 FILLCELL_X16 FILLER_6_318 ();
 FILLCELL_X8 FILLER_6_334 ();
 FILLCELL_X4 FILLER_6_342 ();
 FILLCELL_X1 FILLER_6_346 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X8 FILLER_7_129 ();
 FILLCELL_X2 FILLER_7_137 ();
 FILLCELL_X2 FILLER_7_156 ();
 FILLCELL_X1 FILLER_7_158 ();
 FILLCELL_X8 FILLER_7_170 ();
 FILLCELL_X4 FILLER_7_178 ();
 FILLCELL_X2 FILLER_7_182 ();
 FILLCELL_X2 FILLER_7_201 ();
 FILLCELL_X32 FILLER_7_207 ();
 FILLCELL_X32 FILLER_7_239 ();
 FILLCELL_X8 FILLER_7_271 ();
 FILLCELL_X2 FILLER_7_279 ();
 FILLCELL_X1 FILLER_7_281 ();
 FILLCELL_X32 FILLER_7_299 ();
 FILLCELL_X16 FILLER_7_331 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X16 FILLER_8_129 ();
 FILLCELL_X4 FILLER_8_145 ();
 FILLCELL_X2 FILLER_8_149 ();
 FILLCELL_X1 FILLER_8_151 ();
 FILLCELL_X8 FILLER_8_169 ();
 FILLCELL_X2 FILLER_8_177 ();
 FILLCELL_X1 FILLER_8_179 ();
 FILLCELL_X32 FILLER_8_184 ();
 FILLCELL_X32 FILLER_8_216 ();
 FILLCELL_X32 FILLER_8_248 ();
 FILLCELL_X32 FILLER_8_280 ();
 FILLCELL_X32 FILLER_8_312 ();
 FILLCELL_X2 FILLER_8_344 ();
 FILLCELL_X1 FILLER_8_346 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X16 FILLER_9_129 ();
 FILLCELL_X8 FILLER_9_145 ();
 FILLCELL_X2 FILLER_9_153 ();
 FILLCELL_X32 FILLER_9_163 ();
 FILLCELL_X32 FILLER_9_195 ();
 FILLCELL_X32 FILLER_9_227 ();
 FILLCELL_X8 FILLER_9_259 ();
 FILLCELL_X2 FILLER_9_267 ();
 FILLCELL_X32 FILLER_9_287 ();
 FILLCELL_X2 FILLER_9_319 ();
 FILLCELL_X1 FILLER_9_321 ();
 FILLCELL_X8 FILLER_9_339 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X4 FILLER_10_257 ();
 FILLCELL_X8 FILLER_10_266 ();
 FILLCELL_X4 FILLER_10_291 ();
 FILLCELL_X2 FILLER_10_344 ();
 FILLCELL_X1 FILLER_10_346 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X16 FILLER_11_289 ();
 FILLCELL_X2 FILLER_11_305 ();
 FILLCELL_X1 FILLER_11_307 ();
 FILLCELL_X8 FILLER_11_315 ();
 FILLCELL_X4 FILLER_11_323 ();
 FILLCELL_X2 FILLER_11_327 ();
 FILLCELL_X4 FILLER_11_336 ();
 FILLCELL_X1 FILLER_11_340 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X8 FILLER_12_321 ();
 FILLCELL_X4 FILLER_12_329 ();
 FILLCELL_X2 FILLER_12_333 ();
 FILLCELL_X2 FILLER_12_341 ();
 FILLCELL_X1 FILLER_12_343 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X16 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_145 ();
 FILLCELL_X4 FILLER_13_153 ();
 FILLCELL_X1 FILLER_13_157 ();
 FILLCELL_X32 FILLER_13_162 ();
 FILLCELL_X32 FILLER_13_194 ();
 FILLCELL_X32 FILLER_13_226 ();
 FILLCELL_X32 FILLER_13_258 ();
 FILLCELL_X32 FILLER_13_290 ();
 FILLCELL_X16 FILLER_13_322 ();
 FILLCELL_X8 FILLER_13_338 ();
 FILLCELL_X1 FILLER_13_346 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_161 ();
 FILLCELL_X8 FILLER_14_176 ();
 FILLCELL_X2 FILLER_14_184 ();
 FILLCELL_X32 FILLER_14_199 ();
 FILLCELL_X32 FILLER_14_231 ();
 FILLCELL_X16 FILLER_14_263 ();
 FILLCELL_X8 FILLER_14_279 ();
 FILLCELL_X2 FILLER_14_287 ();
 FILLCELL_X32 FILLER_14_293 ();
 FILLCELL_X16 FILLER_14_325 ();
 FILLCELL_X4 FILLER_14_341 ();
 FILLCELL_X2 FILLER_14_345 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X8 FILLER_15_113 ();
 FILLCELL_X2 FILLER_15_121 ();
 FILLCELL_X1 FILLER_15_123 ();
 FILLCELL_X16 FILLER_15_132 ();
 FILLCELL_X4 FILLER_15_148 ();
 FILLCELL_X2 FILLER_15_152 ();
 FILLCELL_X32 FILLER_15_165 ();
 FILLCELL_X32 FILLER_15_197 ();
 FILLCELL_X32 FILLER_15_229 ();
 FILLCELL_X16 FILLER_15_261 ();
 FILLCELL_X8 FILLER_15_277 ();
 FILLCELL_X1 FILLER_15_285 ();
 FILLCELL_X2 FILLER_15_303 ();
 FILLCELL_X2 FILLER_15_316 ();
 FILLCELL_X1 FILLER_15_318 ();
 FILLCELL_X8 FILLER_15_336 ();
 FILLCELL_X2 FILLER_15_344 ();
 FILLCELL_X1 FILLER_15_346 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X16 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_145 ();
 FILLCELL_X1 FILLER_16_153 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X8 FILLER_16_257 ();
 FILLCELL_X4 FILLER_16_265 ();
 FILLCELL_X2 FILLER_16_269 ();
 FILLCELL_X4 FILLER_16_306 ();
 FILLCELL_X4 FILLER_16_324 ();
 FILLCELL_X1 FILLER_16_328 ();
 FILLCELL_X1 FILLER_16_343 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_17 ();
 FILLCELL_X2 FILLER_17_21 ();
 FILLCELL_X1 FILLER_17_23 ();
 FILLCELL_X32 FILLER_17_41 ();
 FILLCELL_X32 FILLER_17_73 ();
 FILLCELL_X32 FILLER_17_105 ();
 FILLCELL_X32 FILLER_17_137 ();
 FILLCELL_X32 FILLER_17_169 ();
 FILLCELL_X32 FILLER_17_201 ();
 FILLCELL_X32 FILLER_17_233 ();
 FILLCELL_X32 FILLER_17_265 ();
 FILLCELL_X16 FILLER_17_297 ();
 FILLCELL_X4 FILLER_17_313 ();
 FILLCELL_X2 FILLER_17_324 ();
 FILLCELL_X1 FILLER_17_343 ();
 FILLCELL_X2 FILLER_18_7 ();
 FILLCELL_X1 FILLER_18_26 ();
 FILLCELL_X32 FILLER_18_31 ();
 FILLCELL_X32 FILLER_18_63 ();
 FILLCELL_X8 FILLER_18_95 ();
 FILLCELL_X1 FILLER_18_103 ();
 FILLCELL_X2 FILLER_18_115 ();
 FILLCELL_X32 FILLER_18_134 ();
 FILLCELL_X32 FILLER_18_166 ();
 FILLCELL_X32 FILLER_18_198 ();
 FILLCELL_X32 FILLER_18_230 ();
 FILLCELL_X32 FILLER_18_262 ();
 FILLCELL_X16 FILLER_18_294 ();
 FILLCELL_X4 FILLER_18_310 ();
 FILLCELL_X2 FILLER_18_331 ();
 FILLCELL_X2 FILLER_18_342 ();
 FILLCELL_X1 FILLER_19_4 ();
 FILLCELL_X2 FILLER_19_12 ();
 FILLCELL_X1 FILLER_19_21 ();
 FILLCELL_X1 FILLER_19_29 ();
 FILLCELL_X32 FILLER_19_34 ();
 FILLCELL_X32 FILLER_19_66 ();
 FILLCELL_X4 FILLER_19_98 ();
 FILLCELL_X2 FILLER_19_102 ();
 FILLCELL_X1 FILLER_19_104 ();
 FILLCELL_X32 FILLER_19_109 ();
 FILLCELL_X32 FILLER_19_141 ();
 FILLCELL_X32 FILLER_19_173 ();
 FILLCELL_X32 FILLER_19_205 ();
 FILLCELL_X32 FILLER_19_237 ();
 FILLCELL_X32 FILLER_19_269 ();
 FILLCELL_X32 FILLER_19_301 ();
 FILLCELL_X8 FILLER_19_333 ();
 FILLCELL_X4 FILLER_19_341 ();
 FILLCELL_X2 FILLER_19_345 ();
 FILLCELL_X2 FILLER_20_10 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X4 FILLER_20_113 ();
 FILLCELL_X2 FILLER_20_117 ();
 FILLCELL_X32 FILLER_20_132 ();
 FILLCELL_X32 FILLER_20_164 ();
 FILLCELL_X32 FILLER_20_196 ();
 FILLCELL_X32 FILLER_20_228 ();
 FILLCELL_X32 FILLER_20_260 ();
 FILLCELL_X32 FILLER_20_292 ();
 FILLCELL_X16 FILLER_20_324 ();
 FILLCELL_X4 FILLER_20_340 ();
 FILLCELL_X2 FILLER_20_344 ();
 FILLCELL_X1 FILLER_20_346 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_5 ();
 FILLCELL_X2 FILLER_21_12 ();
 FILLCELL_X1 FILLER_21_14 ();
 FILLCELL_X32 FILLER_21_60 ();
 FILLCELL_X32 FILLER_21_92 ();
 FILLCELL_X8 FILLER_21_124 ();
 FILLCELL_X1 FILLER_21_132 ();
 FILLCELL_X32 FILLER_21_140 ();
 FILLCELL_X2 FILLER_21_172 ();
 FILLCELL_X1 FILLER_21_174 ();
 FILLCELL_X32 FILLER_21_179 ();
 FILLCELL_X32 FILLER_21_211 ();
 FILLCELL_X32 FILLER_21_243 ();
 FILLCELL_X32 FILLER_21_275 ();
 FILLCELL_X2 FILLER_21_307 ();
 FILLCELL_X1 FILLER_21_309 ();
 FILLCELL_X16 FILLER_21_331 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_9 ();
 FILLCELL_X32 FILLER_22_24 ();
 FILLCELL_X32 FILLER_22_56 ();
 FILLCELL_X16 FILLER_22_88 ();
 FILLCELL_X8 FILLER_22_104 ();
 FILLCELL_X1 FILLER_22_112 ();
 FILLCELL_X8 FILLER_22_120 ();
 FILLCELL_X2 FILLER_22_128 ();
 FILLCELL_X1 FILLER_22_130 ();
 FILLCELL_X32 FILLER_22_138 ();
 FILLCELL_X32 FILLER_22_170 ();
 FILLCELL_X32 FILLER_22_202 ();
 FILLCELL_X32 FILLER_22_234 ();
 FILLCELL_X32 FILLER_22_266 ();
 FILLCELL_X8 FILLER_22_298 ();
 FILLCELL_X2 FILLER_22_306 ();
 FILLCELL_X1 FILLER_22_308 ();
 FILLCELL_X2 FILLER_22_330 ();
 FILLCELL_X4 FILLER_22_338 ();
 FILLCELL_X2 FILLER_22_342 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_17 ();
 FILLCELL_X8 FILLER_23_22 ();
 FILLCELL_X1 FILLER_23_30 ();
 FILLCELL_X32 FILLER_23_34 ();
 FILLCELL_X16 FILLER_23_66 ();
 FILLCELL_X8 FILLER_23_82 ();
 FILLCELL_X4 FILLER_23_108 ();
 FILLCELL_X32 FILLER_23_126 ();
 FILLCELL_X4 FILLER_23_158 ();
 FILLCELL_X1 FILLER_23_176 ();
 FILLCELL_X32 FILLER_23_197 ();
 FILLCELL_X32 FILLER_23_229 ();
 FILLCELL_X16 FILLER_23_261 ();
 FILLCELL_X2 FILLER_23_277 ();
 FILLCELL_X1 FILLER_23_279 ();
 FILLCELL_X8 FILLER_23_297 ();
 FILLCELL_X2 FILLER_23_305 ();
 FILLCELL_X1 FILLER_23_307 ();
 FILLCELL_X4 FILLER_23_315 ();
 FILLCELL_X2 FILLER_23_319 ();
 FILLCELL_X1 FILLER_23_321 ();
 FILLCELL_X1 FILLER_23_343 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_9 ();
 FILLCELL_X1 FILLER_24_11 ();
 FILLCELL_X16 FILLER_24_15 ();
 FILLCELL_X8 FILLER_24_31 ();
 FILLCELL_X32 FILLER_24_42 ();
 FILLCELL_X8 FILLER_24_74 ();
 FILLCELL_X4 FILLER_24_82 ();
 FILLCELL_X2 FILLER_24_86 ();
 FILLCELL_X32 FILLER_24_126 ();
 FILLCELL_X16 FILLER_24_158 ();
 FILLCELL_X32 FILLER_24_179 ();
 FILLCELL_X32 FILLER_24_211 ();
 FILLCELL_X32 FILLER_24_243 ();
 FILLCELL_X16 FILLER_24_275 ();
 FILLCELL_X1 FILLER_24_291 ();
 FILLCELL_X2 FILLER_24_316 ();
 FILLCELL_X1 FILLER_24_318 ();
 FILLCELL_X4 FILLER_24_339 ();
 FILLCELL_X1 FILLER_24_343 ();
 FILLCELL_X2 FILLER_25_4 ();
 FILLCELL_X2 FILLER_25_9 ();
 FILLCELL_X1 FILLER_25_11 ();
 FILLCELL_X2 FILLER_25_19 ();
 FILLCELL_X4 FILLER_25_25 ();
 FILLCELL_X2 FILLER_25_29 ();
 FILLCELL_X1 FILLER_25_31 ();
 FILLCELL_X4 FILLER_25_39 ();
 FILLCELL_X2 FILLER_25_43 ();
 FILLCELL_X1 FILLER_25_45 ();
 FILLCELL_X32 FILLER_25_50 ();
 FILLCELL_X16 FILLER_25_82 ();
 FILLCELL_X4 FILLER_25_98 ();
 FILLCELL_X2 FILLER_25_102 ();
 FILLCELL_X1 FILLER_25_104 ();
 FILLCELL_X32 FILLER_25_109 ();
 FILLCELL_X32 FILLER_25_141 ();
 FILLCELL_X8 FILLER_25_173 ();
 FILLCELL_X4 FILLER_25_181 ();
 FILLCELL_X32 FILLER_25_189 ();
 FILLCELL_X32 FILLER_25_221 ();
 FILLCELL_X32 FILLER_25_253 ();
 FILLCELL_X1 FILLER_25_285 ();
 FILLCELL_X2 FILLER_25_294 ();
 FILLCELL_X32 FILLER_25_306 ();
 FILLCELL_X8 FILLER_25_338 ();
 FILLCELL_X1 FILLER_25_346 ();
 FILLCELL_X1 FILLER_26_11 ();
 FILLCELL_X8 FILLER_26_39 ();
 FILLCELL_X1 FILLER_26_47 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X16 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_145 ();
 FILLCELL_X32 FILLER_26_157 ();
 FILLCELL_X32 FILLER_26_189 ();
 FILLCELL_X32 FILLER_26_221 ();
 FILLCELL_X32 FILLER_26_253 ();
 FILLCELL_X16 FILLER_26_285 ();
 FILLCELL_X8 FILLER_26_301 ();
 FILLCELL_X4 FILLER_26_309 ();
 FILLCELL_X2 FILLER_26_313 ();
 FILLCELL_X16 FILLER_26_318 ();
 FILLCELL_X8 FILLER_26_334 ();
 FILLCELL_X4 FILLER_26_342 ();
 FILLCELL_X1 FILLER_26_346 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_5 ();
 FILLCELL_X1 FILLER_27_7 ();
 FILLCELL_X4 FILLER_27_11 ();
 FILLCELL_X2 FILLER_27_15 ();
 FILLCELL_X1 FILLER_27_17 ();
 FILLCELL_X32 FILLER_27_21 ();
 FILLCELL_X32 FILLER_27_53 ();
 FILLCELL_X32 FILLER_27_85 ();
 FILLCELL_X32 FILLER_27_117 ();
 FILLCELL_X32 FILLER_27_149 ();
 FILLCELL_X32 FILLER_27_181 ();
 FILLCELL_X32 FILLER_27_213 ();
 FILLCELL_X32 FILLER_27_245 ();
 FILLCELL_X8 FILLER_27_277 ();
 FILLCELL_X2 FILLER_27_285 ();
 FILLCELL_X1 FILLER_27_287 ();
 FILLCELL_X2 FILLER_27_327 ();
 FILLCELL_X2 FILLER_27_342 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_5 ();
 FILLCELL_X1 FILLER_28_26 ();
 FILLCELL_X4 FILLER_28_34 ();
 FILLCELL_X1 FILLER_28_38 ();
 FILLCELL_X32 FILLER_28_43 ();
 FILLCELL_X32 FILLER_28_75 ();
 FILLCELL_X32 FILLER_28_107 ();
 FILLCELL_X32 FILLER_28_139 ();
 FILLCELL_X32 FILLER_28_171 ();
 FILLCELL_X32 FILLER_28_203 ();
 FILLCELL_X32 FILLER_28_235 ();
 FILLCELL_X32 FILLER_28_267 ();
 FILLCELL_X16 FILLER_28_299 ();
 FILLCELL_X2 FILLER_28_315 ();
 FILLCELL_X4 FILLER_28_341 ();
 FILLCELL_X2 FILLER_28_345 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_9 ();
 FILLCELL_X16 FILLER_29_21 ();
 FILLCELL_X1 FILLER_29_37 ();
 FILLCELL_X32 FILLER_29_55 ();
 FILLCELL_X32 FILLER_29_87 ();
 FILLCELL_X32 FILLER_29_119 ();
 FILLCELL_X32 FILLER_29_151 ();
 FILLCELL_X32 FILLER_29_183 ();
 FILLCELL_X32 FILLER_29_215 ();
 FILLCELL_X32 FILLER_29_247 ();
 FILLCELL_X32 FILLER_29_279 ();
 FILLCELL_X16 FILLER_29_311 ();
 FILLCELL_X1 FILLER_29_327 ();
 FILLCELL_X4 FILLER_29_331 ();
 FILLCELL_X2 FILLER_29_335 ();
 FILLCELL_X1 FILLER_29_337 ();
 FILLCELL_X2 FILLER_29_344 ();
 FILLCELL_X1 FILLER_29_346 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X4 FILLER_30_9 ();
 FILLCELL_X2 FILLER_30_13 ();
 FILLCELL_X32 FILLER_30_32 ();
 FILLCELL_X32 FILLER_30_64 ();
 FILLCELL_X32 FILLER_30_96 ();
 FILLCELL_X32 FILLER_30_128 ();
 FILLCELL_X32 FILLER_30_160 ();
 FILLCELL_X32 FILLER_30_192 ();
 FILLCELL_X32 FILLER_30_224 ();
 FILLCELL_X32 FILLER_30_256 ();
 FILLCELL_X2 FILLER_30_288 ();
 FILLCELL_X8 FILLER_30_294 ();
 FILLCELL_X1 FILLER_30_302 ();
 FILLCELL_X4 FILLER_30_310 ();
 FILLCELL_X2 FILLER_30_314 ();
 FILLCELL_X2 FILLER_30_327 ();
 FILLCELL_X1 FILLER_30_343 ();
 FILLCELL_X1 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_5 ();
 FILLCELL_X32 FILLER_31_37 ();
 FILLCELL_X32 FILLER_31_69 ();
 FILLCELL_X32 FILLER_31_101 ();
 FILLCELL_X32 FILLER_31_133 ();
 FILLCELL_X32 FILLER_31_165 ();
 FILLCELL_X32 FILLER_31_197 ();
 FILLCELL_X32 FILLER_31_229 ();
 FILLCELL_X16 FILLER_31_261 ();
 FILLCELL_X8 FILLER_31_277 ();
 FILLCELL_X1 FILLER_31_285 ();
 FILLCELL_X8 FILLER_31_303 ();
 FILLCELL_X4 FILLER_31_311 ();
 FILLCELL_X2 FILLER_31_315 ();
 FILLCELL_X1 FILLER_31_317 ();
 FILLCELL_X8 FILLER_31_335 ();
 FILLCELL_X4 FILLER_31_343 ();
 FILLCELL_X2 FILLER_32_4 ();
 FILLCELL_X1 FILLER_32_6 ();
 FILLCELL_X2 FILLER_32_10 ();
 FILLCELL_X32 FILLER_32_19 ();
 FILLCELL_X32 FILLER_32_51 ();
 FILLCELL_X32 FILLER_32_83 ();
 FILLCELL_X32 FILLER_32_115 ();
 FILLCELL_X32 FILLER_32_147 ();
 FILLCELL_X32 FILLER_32_179 ();
 FILLCELL_X32 FILLER_32_211 ();
 FILLCELL_X32 FILLER_32_243 ();
 FILLCELL_X32 FILLER_32_275 ();
 FILLCELL_X32 FILLER_32_307 ();
 FILLCELL_X8 FILLER_32_339 ();
 FILLCELL_X2 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_3 ();
 FILLCELL_X32 FILLER_33_31 ();
 FILLCELL_X16 FILLER_33_63 ();
 FILLCELL_X8 FILLER_33_79 ();
 FILLCELL_X2 FILLER_33_87 ();
 FILLCELL_X32 FILLER_33_96 ();
 FILLCELL_X32 FILLER_33_128 ();
 FILLCELL_X32 FILLER_33_160 ();
 FILLCELL_X32 FILLER_33_192 ();
 FILLCELL_X32 FILLER_33_224 ();
 FILLCELL_X32 FILLER_33_256 ();
 FILLCELL_X32 FILLER_33_288 ();
 FILLCELL_X16 FILLER_33_320 ();
 FILLCELL_X1 FILLER_33_336 ();
 FILLCELL_X4 FILLER_33_340 ();
 FILLCELL_X2 FILLER_33_344 ();
 FILLCELL_X1 FILLER_33_346 ();
 FILLCELL_X8 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_9 ();
 FILLCELL_X32 FILLER_34_29 ();
 FILLCELL_X32 FILLER_34_61 ();
 FILLCELL_X32 FILLER_34_93 ();
 FILLCELL_X32 FILLER_34_125 ();
 FILLCELL_X32 FILLER_34_157 ();
 FILLCELL_X32 FILLER_34_189 ();
 FILLCELL_X32 FILLER_34_221 ();
 FILLCELL_X32 FILLER_34_253 ();
 FILLCELL_X16 FILLER_34_285 ();
 FILLCELL_X8 FILLER_34_301 ();
 FILLCELL_X4 FILLER_34_309 ();
 FILLCELL_X1 FILLER_34_313 ();
 FILLCELL_X4 FILLER_34_325 ();
 FILLCELL_X2 FILLER_34_336 ();
 FILLCELL_X1 FILLER_34_338 ();
 FILLCELL_X2 FILLER_34_342 ();
 FILLCELL_X8 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_9 ();
 FILLCELL_X32 FILLER_35_31 ();
 FILLCELL_X32 FILLER_35_63 ();
 FILLCELL_X32 FILLER_35_95 ();
 FILLCELL_X32 FILLER_35_127 ();
 FILLCELL_X32 FILLER_35_159 ();
 FILLCELL_X32 FILLER_35_191 ();
 FILLCELL_X16 FILLER_35_223 ();
 FILLCELL_X8 FILLER_35_239 ();
 FILLCELL_X1 FILLER_35_247 ();
 FILLCELL_X32 FILLER_35_256 ();
 FILLCELL_X16 FILLER_35_288 ();
 FILLCELL_X8 FILLER_35_304 ();
 FILLCELL_X4 FILLER_35_312 ();
 FILLCELL_X2 FILLER_35_316 ();
 FILLCELL_X1 FILLER_35_318 ();
 FILLCELL_X4 FILLER_35_343 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X16 FILLER_36_321 ();
 FILLCELL_X8 FILLER_36_337 ();
 FILLCELL_X2 FILLER_36_345 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X16 FILLER_37_193 ();
 FILLCELL_X8 FILLER_37_209 ();
 FILLCELL_X2 FILLER_37_217 ();
 FILLCELL_X1 FILLER_37_219 ();
 FILLCELL_X32 FILLER_37_224 ();
 FILLCELL_X32 FILLER_37_256 ();
 FILLCELL_X32 FILLER_37_288 ();
 FILLCELL_X16 FILLER_37_320 ();
 FILLCELL_X8 FILLER_37_336 ();
 FILLCELL_X2 FILLER_37_344 ();
 FILLCELL_X1 FILLER_37_346 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_20 ();
 FILLCELL_X32 FILLER_38_52 ();
 FILLCELL_X4 FILLER_38_84 ();
 FILLCELL_X2 FILLER_38_88 ();
 FILLCELL_X1 FILLER_38_90 ();
 FILLCELL_X32 FILLER_38_125 ();
 FILLCELL_X16 FILLER_38_157 ();
 FILLCELL_X8 FILLER_38_173 ();
 FILLCELL_X1 FILLER_38_181 ();
 FILLCELL_X8 FILLER_38_203 ();
 FILLCELL_X4 FILLER_38_211 ();
 FILLCELL_X1 FILLER_38_215 ();
 FILLCELL_X32 FILLER_38_233 ();
 FILLCELL_X32 FILLER_38_265 ();
 FILLCELL_X32 FILLER_38_297 ();
 FILLCELL_X16 FILLER_38_329 ();
 FILLCELL_X2 FILLER_38_345 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_17 ();
 FILLCELL_X1 FILLER_39_19 ();
 FILLCELL_X32 FILLER_39_27 ();
 FILLCELL_X32 FILLER_39_59 ();
 FILLCELL_X4 FILLER_39_91 ();
 FILLCELL_X1 FILLER_39_95 ();
 FILLCELL_X1 FILLER_39_100 ();
 FILLCELL_X2 FILLER_39_110 ();
 FILLCELL_X1 FILLER_39_112 ();
 FILLCELL_X8 FILLER_39_120 ();
 FILLCELL_X2 FILLER_39_128 ();
 FILLCELL_X4 FILLER_39_144 ();
 FILLCELL_X1 FILLER_39_148 ();
 FILLCELL_X16 FILLER_39_153 ();
 FILLCELL_X8 FILLER_39_169 ();
 FILLCELL_X8 FILLER_39_184 ();
 FILLCELL_X8 FILLER_39_213 ();
 FILLCELL_X2 FILLER_39_233 ();
 FILLCELL_X8 FILLER_39_252 ();
 FILLCELL_X4 FILLER_39_260 ();
 FILLCELL_X1 FILLER_39_264 ();
 FILLCELL_X8 FILLER_39_269 ();
 FILLCELL_X4 FILLER_39_277 ();
 FILLCELL_X2 FILLER_39_281 ();
 FILLCELL_X32 FILLER_39_311 ();
 FILLCELL_X4 FILLER_39_343 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X8 FILLER_40_17 ();
 FILLCELL_X32 FILLER_40_29 ();
 FILLCELL_X32 FILLER_40_61 ();
 FILLCELL_X8 FILLER_40_93 ();
 FILLCELL_X2 FILLER_40_101 ();
 FILLCELL_X1 FILLER_40_103 ();
 FILLCELL_X32 FILLER_40_115 ();
 FILLCELL_X1 FILLER_40_147 ();
 FILLCELL_X16 FILLER_40_165 ();
 FILLCELL_X4 FILLER_40_181 ();
 FILLCELL_X2 FILLER_40_185 ();
 FILLCELL_X1 FILLER_40_187 ();
 FILLCELL_X16 FILLER_40_195 ();
 FILLCELL_X4 FILLER_40_211 ();
 FILLCELL_X2 FILLER_40_222 ();
 FILLCELL_X1 FILLER_40_224 ();
 FILLCELL_X16 FILLER_40_232 ();
 FILLCELL_X8 FILLER_40_248 ();
 FILLCELL_X4 FILLER_40_256 ();
 FILLCELL_X2 FILLER_40_260 ();
 FILLCELL_X32 FILLER_40_279 ();
 FILLCELL_X32 FILLER_40_311 ();
 FILLCELL_X4 FILLER_40_343 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X4 FILLER_41_17 ();
 FILLCELL_X1 FILLER_41_21 ();
 FILLCELL_X16 FILLER_41_39 ();
 FILLCELL_X8 FILLER_41_55 ();
 FILLCELL_X4 FILLER_41_63 ();
 FILLCELL_X2 FILLER_41_67 ();
 FILLCELL_X8 FILLER_41_90 ();
 FILLCELL_X4 FILLER_41_98 ();
 FILLCELL_X32 FILLER_41_119 ();
 FILLCELL_X32 FILLER_41_151 ();
 FILLCELL_X32 FILLER_41_183 ();
 FILLCELL_X32 FILLER_41_215 ();
 FILLCELL_X16 FILLER_41_247 ();
 FILLCELL_X32 FILLER_41_270 ();
 FILLCELL_X32 FILLER_41_302 ();
 FILLCELL_X8 FILLER_41_334 ();
 FILLCELL_X4 FILLER_41_342 ();
 FILLCELL_X1 FILLER_41_346 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X16 FILLER_42_65 ();
 FILLCELL_X2 FILLER_42_81 ();
 FILLCELL_X16 FILLER_42_90 ();
 FILLCELL_X8 FILLER_42_106 ();
 FILLCELL_X2 FILLER_42_114 ();
 FILLCELL_X1 FILLER_42_116 ();
 FILLCELL_X32 FILLER_42_124 ();
 FILLCELL_X16 FILLER_42_156 ();
 FILLCELL_X4 FILLER_42_172 ();
 FILLCELL_X2 FILLER_42_176 ();
 FILLCELL_X1 FILLER_42_178 ();
 FILLCELL_X4 FILLER_42_194 ();
 FILLCELL_X16 FILLER_42_205 ();
 FILLCELL_X4 FILLER_42_221 ();
 FILLCELL_X32 FILLER_42_236 ();
 FILLCELL_X32 FILLER_42_268 ();
 FILLCELL_X32 FILLER_42_300 ();
 FILLCELL_X8 FILLER_42_332 ();
 FILLCELL_X4 FILLER_42_340 ();
 FILLCELL_X2 FILLER_42_344 ();
 FILLCELL_X1 FILLER_42_346 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X8 FILLER_43_33 ();
 FILLCELL_X2 FILLER_43_41 ();
 FILLCELL_X32 FILLER_43_47 ();
 FILLCELL_X16 FILLER_43_79 ();
 FILLCELL_X8 FILLER_43_95 ();
 FILLCELL_X4 FILLER_43_103 ();
 FILLCELL_X2 FILLER_43_107 ();
 FILLCELL_X8 FILLER_43_113 ();
 FILLCELL_X4 FILLER_43_121 ();
 FILLCELL_X4 FILLER_43_132 ();
 FILLCELL_X2 FILLER_43_136 ();
 FILLCELL_X16 FILLER_43_149 ();
 FILLCELL_X4 FILLER_43_165 ();
 FILLCELL_X16 FILLER_43_203 ();
 FILLCELL_X2 FILLER_43_219 ();
 FILLCELL_X1 FILLER_43_221 ();
 FILLCELL_X1 FILLER_43_246 ();
 FILLCELL_X32 FILLER_43_251 ();
 FILLCELL_X32 FILLER_43_283 ();
 FILLCELL_X32 FILLER_43_315 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X4 FILLER_44_33 ();
 FILLCELL_X16 FILLER_44_68 ();
 FILLCELL_X4 FILLER_44_102 ();
 FILLCELL_X1 FILLER_44_106 ();
 FILLCELL_X4 FILLER_44_124 ();
 FILLCELL_X16 FILLER_44_159 ();
 FILLCELL_X2 FILLER_44_175 ();
 FILLCELL_X1 FILLER_44_177 ();
 FILLCELL_X4 FILLER_44_185 ();
 FILLCELL_X2 FILLER_44_189 ();
 FILLCELL_X1 FILLER_44_191 ();
 FILLCELL_X16 FILLER_44_206 ();
 FILLCELL_X2 FILLER_44_243 ();
 FILLCELL_X1 FILLER_44_245 ();
 FILLCELL_X2 FILLER_44_263 ();
 FILLCELL_X1 FILLER_44_265 ();
 FILLCELL_X1 FILLER_44_273 ();
 FILLCELL_X32 FILLER_44_285 ();
 FILLCELL_X16 FILLER_44_317 ();
 FILLCELL_X8 FILLER_44_333 ();
 FILLCELL_X4 FILLER_44_341 ();
 FILLCELL_X2 FILLER_44_345 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X16 FILLER_45_33 ();
 FILLCELL_X4 FILLER_45_49 ();
 FILLCELL_X2 FILLER_45_53 ();
 FILLCELL_X1 FILLER_45_55 ();
 FILLCELL_X16 FILLER_45_63 ();
 FILLCELL_X4 FILLER_45_79 ();
 FILLCELL_X2 FILLER_45_83 ();
 FILLCELL_X4 FILLER_45_92 ();
 FILLCELL_X8 FILLER_45_113 ();
 FILLCELL_X4 FILLER_45_121 ();
 FILLCELL_X1 FILLER_45_132 ();
 FILLCELL_X32 FILLER_45_147 ();
 FILLCELL_X2 FILLER_45_179 ();
 FILLCELL_X1 FILLER_45_181 ();
 FILLCELL_X16 FILLER_45_195 ();
 FILLCELL_X8 FILLER_45_211 ();
 FILLCELL_X4 FILLER_45_219 ();
 FILLCELL_X2 FILLER_45_226 ();
 FILLCELL_X1 FILLER_45_231 ();
 FILLCELL_X16 FILLER_45_239 ();
 FILLCELL_X8 FILLER_45_255 ();
 FILLCELL_X4 FILLER_45_263 ();
 FILLCELL_X2 FILLER_45_267 ();
 FILLCELL_X1 FILLER_45_269 ();
 FILLCELL_X32 FILLER_45_294 ();
 FILLCELL_X16 FILLER_45_326 ();
 FILLCELL_X4 FILLER_45_342 ();
 FILLCELL_X1 FILLER_45_346 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X16 FILLER_46_33 ();
 FILLCELL_X8 FILLER_46_49 ();
 FILLCELL_X2 FILLER_46_57 ();
 FILLCELL_X16 FILLER_46_68 ();
 FILLCELL_X4 FILLER_46_84 ();
 FILLCELL_X2 FILLER_46_88 ();
 FILLCELL_X2 FILLER_46_96 ();
 FILLCELL_X1 FILLER_46_98 ();
 FILLCELL_X4 FILLER_46_102 ();
 FILLCELL_X2 FILLER_46_109 ();
 FILLCELL_X2 FILLER_46_114 ();
 FILLCELL_X4 FILLER_46_122 ();
 FILLCELL_X2 FILLER_46_126 ();
 FILLCELL_X1 FILLER_46_128 ();
 FILLCELL_X1 FILLER_46_141 ();
 FILLCELL_X2 FILLER_46_145 ();
 FILLCELL_X1 FILLER_46_150 ();
 FILLCELL_X16 FILLER_46_160 ();
 FILLCELL_X2 FILLER_46_176 ();
 FILLCELL_X1 FILLER_46_181 ();
 FILLCELL_X2 FILLER_46_191 ();
 FILLCELL_X16 FILLER_46_199 ();
 FILLCELL_X1 FILLER_46_215 ();
 FILLCELL_X4 FILLER_46_219 ();
 FILLCELL_X2 FILLER_46_229 ();
 FILLCELL_X4 FILLER_46_237 ();
 FILLCELL_X16 FILLER_46_244 ();
 FILLCELL_X1 FILLER_46_260 ();
 FILLCELL_X2 FILLER_46_267 ();
 FILLCELL_X32 FILLER_46_278 ();
 FILLCELL_X32 FILLER_46_310 ();
 FILLCELL_X4 FILLER_46_342 ();
 FILLCELL_X1 FILLER_46_346 ();
endmodule
