module bidirectional_shift_register (clk,
    direction,
    enable,
    load_en,
    rst_n,
    serial_in,
    shift_en,
    parallel_in,
    parallel_out);
 input clk;
 input direction;
 input enable;
 input load_en;
 input rst_n;
 input serial_in;
 input shift_en;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _057_ (.A(rst_n),
    .Z(_008_));
 BUF_X4 _058_ (.A(net2),
    .Z(_009_));
 OAI21_X4 _059_ (.A(net1),
    .B1(_009_),
    .B2(net12),
    .ZN(_010_));
 NAND3_X1 _060_ (.A1(net13),
    .A2(_008_),
    .A3(_010_),
    .ZN(_011_));
 BUF_X2 _061_ (.A(direction),
    .Z(_012_));
 MUX2_X1 _062_ (.A(net14),
    .B(net11),
    .S(_012_),
    .Z(_013_));
 NOR2_X1 _063_ (.A1(_009_),
    .A2(_013_),
    .ZN(_014_));
 OR2_X1 _064_ (.A1(net12),
    .A2(net2),
    .ZN(_015_));
 BUF_X4 _065_ (.A(_015_),
    .Z(_016_));
 AND2_X2 _066_ (.A1(net1),
    .A2(_008_),
    .ZN(_017_));
 BUF_X16 _067_ (.A(_017_),
    .Z(_018_));
 INV_X4 _068_ (.A(_009_),
    .ZN(_019_));
 OAI211_X2 _069_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net3),
    .ZN(_020_));
 OAI21_X1 _070_ (.A(_011_),
    .B1(_014_),
    .B2(_020_),
    .ZN(_000_));
 NAND3_X1 _071_ (.A1(net14),
    .A2(_008_),
    .A3(_010_),
    .ZN(_021_));
 MUX2_X1 _072_ (.A(net15),
    .B(net13),
    .S(_012_),
    .Z(_022_));
 NOR2_X1 _073_ (.A1(_009_),
    .A2(_022_),
    .ZN(_023_));
 OAI211_X2 _074_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net4),
    .ZN(_024_));
 OAI21_X1 _075_ (.A(_021_),
    .B1(_023_),
    .B2(_024_),
    .ZN(_001_));
 NAND3_X1 _076_ (.A1(net15),
    .A2(_008_),
    .A3(_010_),
    .ZN(_025_));
 MUX2_X1 _077_ (.A(net16),
    .B(net14),
    .S(_012_),
    .Z(_026_));
 NOR2_X1 _078_ (.A1(_009_),
    .A2(_026_),
    .ZN(_027_));
 OAI211_X2 _079_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net5),
    .ZN(_028_));
 OAI21_X1 _080_ (.A(_025_),
    .B1(_027_),
    .B2(_028_),
    .ZN(_002_));
 NAND3_X1 _081_ (.A1(net16),
    .A2(_008_),
    .A3(_010_),
    .ZN(_029_));
 MUX2_X1 _082_ (.A(net17),
    .B(net15),
    .S(_012_),
    .Z(_030_));
 NOR2_X1 _083_ (.A1(_009_),
    .A2(_030_),
    .ZN(_031_));
 OAI211_X2 _084_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net6),
    .ZN(_032_));
 OAI21_X1 _085_ (.A(_029_),
    .B1(_031_),
    .B2(_032_),
    .ZN(_003_));
 NAND3_X1 _086_ (.A1(net17),
    .A2(_008_),
    .A3(_010_),
    .ZN(_033_));
 MUX2_X1 _087_ (.A(net18),
    .B(net16),
    .S(_012_),
    .Z(_034_));
 NOR2_X1 _088_ (.A1(_009_),
    .A2(_034_),
    .ZN(_035_));
 OAI211_X2 _089_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net7),
    .ZN(_036_));
 OAI21_X1 _090_ (.A(_033_),
    .B1(_035_),
    .B2(_036_),
    .ZN(_004_));
 NAND3_X1 _091_ (.A1(net18),
    .A2(_008_),
    .A3(_010_),
    .ZN(_037_));
 MUX2_X1 _092_ (.A(net19),
    .B(net17),
    .S(_012_),
    .Z(_038_));
 NOR2_X1 _093_ (.A1(_009_),
    .A2(_038_),
    .ZN(_039_));
 OAI211_X2 _094_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net8),
    .ZN(_040_));
 OAI21_X1 _095_ (.A(_037_),
    .B1(_039_),
    .B2(_040_),
    .ZN(_005_));
 NAND3_X1 _096_ (.A1(net19),
    .A2(_008_),
    .A3(_010_),
    .ZN(_041_));
 MUX2_X1 _097_ (.A(net20),
    .B(net18),
    .S(_012_),
    .Z(_042_));
 NOR2_X1 _098_ (.A1(_009_),
    .A2(_042_),
    .ZN(_043_));
 OAI211_X2 _099_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net9),
    .ZN(_044_));
 OAI21_X1 _100_ (.A(_041_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_006_));
 NAND3_X1 _101_ (.A1(net20),
    .A2(_008_),
    .A3(_010_),
    .ZN(_045_));
 MUX2_X1 _102_ (.A(net11),
    .B(net19),
    .S(_012_),
    .Z(_046_));
 NOR2_X1 _103_ (.A1(_009_),
    .A2(_046_),
    .ZN(_047_));
 OAI211_X2 _104_ (.A(_016_),
    .B(_018_),
    .C1(_019_),
    .C2(net10),
    .ZN(_048_));
 OAI21_X1 _105_ (.A(_045_),
    .B1(_047_),
    .B2(_048_),
    .ZN(_007_));
 DFF_X1 \parallel_out[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_056_));
 DFF_X1 \parallel_out[1]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_055_));
 DFF_X1 \parallel_out[2]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_054_));
 DFF_X1 \parallel_out[3]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_053_));
 DFF_X1 \parallel_out[4]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_052_));
 DFF_X1 \parallel_out[5]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net18),
    .QN(_051_));
 DFF_X1 \parallel_out[6]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_050_));
 DFF_X1 \parallel_out[7]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net20),
    .QN(_049_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_67 ();
 BUF_X1 input1 (.A(enable),
    .Z(net1));
 BUF_X1 input2 (.A(load_en),
    .Z(net2));
 BUF_X1 input3 (.A(parallel_in[0]),
    .Z(net3));
 BUF_X1 input4 (.A(parallel_in[1]),
    .Z(net4));
 BUF_X1 input5 (.A(parallel_in[2]),
    .Z(net5));
 BUF_X1 input6 (.A(parallel_in[3]),
    .Z(net6));
 BUF_X1 input7 (.A(parallel_in[4]),
    .Z(net7));
 BUF_X1 input8 (.A(parallel_in[5]),
    .Z(net8));
 BUF_X1 input9 (.A(parallel_in[6]),
    .Z(net9));
 BUF_X1 input10 (.A(parallel_in[7]),
    .Z(net10));
 BUF_X1 input11 (.A(serial_in),
    .Z(net11));
 BUF_X1 input12 (.A(shift_en),
    .Z(net12));
 BUF_X1 output13 (.A(net13),
    .Z(parallel_out[0]));
 BUF_X1 output14 (.A(net14),
    .Z(parallel_out[1]));
 BUF_X1 output15 (.A(net15),
    .Z(parallel_out[2]));
 BUF_X1 output16 (.A(net16),
    .Z(parallel_out[3]));
 BUF_X1 output17 (.A(net17),
    .Z(parallel_out[4]));
 BUF_X1 output18 (.A(net18),
    .Z(parallel_out[5]));
 BUF_X1 output19 (.A(net19),
    .Z(parallel_out[6]));
 BUF_X1 output20 (.A(net20),
    .Z(parallel_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_113 ();
 FILLCELL_X8 FILLER_0_120 ();
 FILLCELL_X4 FILLER_0_134 ();
 FILLCELL_X1 FILLER_0_141 ();
 FILLCELL_X32 FILLER_0_145 ();
 FILLCELL_X32 FILLER_0_177 ();
 FILLCELL_X32 FILLER_0_209 ();
 FILLCELL_X8 FILLER_0_241 ();
 FILLCELL_X4 FILLER_0_249 ();
 FILLCELL_X2 FILLER_0_253 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X8 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_137 ();
 FILLCELL_X32 FILLER_1_144 ();
 FILLCELL_X32 FILLER_1_176 ();
 FILLCELL_X32 FILLER_1_208 ();
 FILLCELL_X8 FILLER_1_240 ();
 FILLCELL_X4 FILLER_1_248 ();
 FILLCELL_X2 FILLER_1_252 ();
 FILLCELL_X1 FILLER_1_254 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X16 FILLER_2_225 ();
 FILLCELL_X8 FILLER_2_241 ();
 FILLCELL_X4 FILLER_2_249 ();
 FILLCELL_X2 FILLER_2_253 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X16 FILLER_3_225 ();
 FILLCELL_X8 FILLER_3_241 ();
 FILLCELL_X4 FILLER_3_249 ();
 FILLCELL_X2 FILLER_3_253 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X16 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_241 ();
 FILLCELL_X4 FILLER_4_249 ();
 FILLCELL_X2 FILLER_4_253 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X16 FILLER_5_225 ();
 FILLCELL_X8 FILLER_5_241 ();
 FILLCELL_X4 FILLER_5_249 ();
 FILLCELL_X2 FILLER_5_253 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X16 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_241 ();
 FILLCELL_X4 FILLER_6_249 ();
 FILLCELL_X2 FILLER_6_253 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X16 FILLER_7_225 ();
 FILLCELL_X8 FILLER_7_241 ();
 FILLCELL_X4 FILLER_7_249 ();
 FILLCELL_X2 FILLER_7_253 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X8 FILLER_8_97 ();
 FILLCELL_X4 FILLER_8_105 ();
 FILLCELL_X2 FILLER_8_109 ();
 FILLCELL_X32 FILLER_8_118 ();
 FILLCELL_X32 FILLER_8_150 ();
 FILLCELL_X32 FILLER_8_182 ();
 FILLCELL_X32 FILLER_8_214 ();
 FILLCELL_X8 FILLER_8_246 ();
 FILLCELL_X1 FILLER_8_254 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X4 FILLER_9_129 ();
 FILLCELL_X2 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_135 ();
 FILLCELL_X32 FILLER_9_147 ();
 FILLCELL_X32 FILLER_9_179 ();
 FILLCELL_X32 FILLER_9_211 ();
 FILLCELL_X8 FILLER_9_243 ();
 FILLCELL_X4 FILLER_9_251 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X4 FILLER_10_129 ();
 FILLCELL_X2 FILLER_10_133 ();
 FILLCELL_X1 FILLER_10_135 ();
 FILLCELL_X32 FILLER_10_154 ();
 FILLCELL_X32 FILLER_10_186 ();
 FILLCELL_X32 FILLER_10_218 ();
 FILLCELL_X4 FILLER_10_250 ();
 FILLCELL_X1 FILLER_10_254 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_137 ();
 FILLCELL_X8 FILLER_11_148 ();
 FILLCELL_X2 FILLER_11_156 ();
 FILLCELL_X32 FILLER_11_183 ();
 FILLCELL_X32 FILLER_11_215 ();
 FILLCELL_X8 FILLER_11_247 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X2 FILLER_12_121 ();
 FILLCELL_X1 FILLER_12_123 ();
 FILLCELL_X32 FILLER_12_138 ();
 FILLCELL_X32 FILLER_12_170 ();
 FILLCELL_X32 FILLER_12_202 ();
 FILLCELL_X16 FILLER_12_234 ();
 FILLCELL_X4 FILLER_12_250 ();
 FILLCELL_X1 FILLER_12_254 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_124 ();
 FILLCELL_X32 FILLER_13_134 ();
 FILLCELL_X32 FILLER_13_166 ();
 FILLCELL_X32 FILLER_13_198 ();
 FILLCELL_X16 FILLER_13_230 ();
 FILLCELL_X8 FILLER_13_246 ();
 FILLCELL_X1 FILLER_13_254 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_17 ();
 FILLCELL_X32 FILLER_14_28 ();
 FILLCELL_X32 FILLER_14_60 ();
 FILLCELL_X8 FILLER_14_92 ();
 FILLCELL_X16 FILLER_14_121 ();
 FILLCELL_X8 FILLER_14_137 ();
 FILLCELL_X1 FILLER_14_145 ();
 FILLCELL_X2 FILLER_14_154 ();
 FILLCELL_X1 FILLER_14_156 ();
 FILLCELL_X32 FILLER_14_166 ();
 FILLCELL_X16 FILLER_14_198 ();
 FILLCELL_X8 FILLER_14_214 ();
 FILLCELL_X2 FILLER_14_222 ();
 FILLCELL_X1 FILLER_14_224 ();
 FILLCELL_X2 FILLER_14_228 ();
 FILLCELL_X16 FILLER_14_233 ();
 FILLCELL_X4 FILLER_14_249 ();
 FILLCELL_X2 FILLER_14_253 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X1 FILLER_15_117 ();
 FILLCELL_X16 FILLER_15_125 ();
 FILLCELL_X4 FILLER_15_141 ();
 FILLCELL_X2 FILLER_15_145 ();
 FILLCELL_X4 FILLER_15_157 ();
 FILLCELL_X2 FILLER_15_161 ();
 FILLCELL_X1 FILLER_15_163 ();
 FILLCELL_X32 FILLER_15_181 ();
 FILLCELL_X8 FILLER_15_213 ();
 FILLCELL_X4 FILLER_15_221 ();
 FILLCELL_X2 FILLER_15_225 ();
 FILLCELL_X16 FILLER_15_230 ();
 FILLCELL_X8 FILLER_15_246 ();
 FILLCELL_X1 FILLER_15_254 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_97 ();
 FILLCELL_X4 FILLER_16_105 ();
 FILLCELL_X1 FILLER_16_109 ();
 FILLCELL_X1 FILLER_16_117 ();
 FILLCELL_X8 FILLER_16_129 ();
 FILLCELL_X4 FILLER_16_137 ();
 FILLCELL_X2 FILLER_16_141 ();
 FILLCELL_X1 FILLER_16_143 ();
 FILLCELL_X2 FILLER_16_151 ();
 FILLCELL_X1 FILLER_16_153 ();
 FILLCELL_X32 FILLER_16_166 ();
 FILLCELL_X32 FILLER_16_198 ();
 FILLCELL_X16 FILLER_16_230 ();
 FILLCELL_X8 FILLER_16_246 ();
 FILLCELL_X1 FILLER_16_254 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_9 ();
 FILLCELL_X32 FILLER_17_16 ();
 FILLCELL_X32 FILLER_17_48 ();
 FILLCELL_X32 FILLER_17_80 ();
 FILLCELL_X2 FILLER_17_112 ();
 FILLCELL_X16 FILLER_17_131 ();
 FILLCELL_X2 FILLER_17_147 ();
 FILLCELL_X1 FILLER_17_149 ();
 FILLCELL_X1 FILLER_17_154 ();
 FILLCELL_X32 FILLER_17_159 ();
 FILLCELL_X16 FILLER_17_191 ();
 FILLCELL_X8 FILLER_17_207 ();
 FILLCELL_X1 FILLER_17_215 ();
 FILLCELL_X32 FILLER_17_219 ();
 FILLCELL_X4 FILLER_17_251 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_123 ();
 FILLCELL_X8 FILLER_18_155 ();
 FILLCELL_X4 FILLER_18_163 ();
 FILLCELL_X1 FILLER_18_167 ();
 FILLCELL_X16 FILLER_18_190 ();
 FILLCELL_X8 FILLER_18_206 ();
 FILLCELL_X2 FILLER_18_214 ();
 FILLCELL_X32 FILLER_18_219 ();
 FILLCELL_X4 FILLER_18_251 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X16 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_81 ();
 FILLCELL_X4 FILLER_19_89 ();
 FILLCELL_X1 FILLER_19_93 ();
 FILLCELL_X4 FILLER_19_111 ();
 FILLCELL_X16 FILLER_19_123 ();
 FILLCELL_X1 FILLER_19_139 ();
 FILLCELL_X2 FILLER_19_155 ();
 FILLCELL_X32 FILLER_19_166 ();
 FILLCELL_X32 FILLER_19_198 ();
 FILLCELL_X16 FILLER_19_230 ();
 FILLCELL_X8 FILLER_19_246 ();
 FILLCELL_X1 FILLER_19_254 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_5 ();
 FILLCELL_X32 FILLER_20_9 ();
 FILLCELL_X32 FILLER_20_41 ();
 FILLCELL_X32 FILLER_20_73 ();
 FILLCELL_X4 FILLER_20_105 ();
 FILLCELL_X1 FILLER_20_109 ();
 FILLCELL_X1 FILLER_20_126 ();
 FILLCELL_X8 FILLER_20_136 ();
 FILLCELL_X2 FILLER_20_144 ();
 FILLCELL_X1 FILLER_20_150 ();
 FILLCELL_X4 FILLER_20_155 ();
 FILLCELL_X32 FILLER_20_163 ();
 FILLCELL_X32 FILLER_20_195 ();
 FILLCELL_X16 FILLER_20_227 ();
 FILLCELL_X8 FILLER_20_243 ();
 FILLCELL_X4 FILLER_20_251 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_97 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X2 FILLER_21_117 ();
 FILLCELL_X16 FILLER_21_122 ();
 FILLCELL_X4 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_142 ();
 FILLCELL_X8 FILLER_21_146 ();
 FILLCELL_X4 FILLER_21_154 ();
 FILLCELL_X2 FILLER_21_158 ();
 FILLCELL_X1 FILLER_21_160 ();
 FILLCELL_X32 FILLER_21_178 ();
 FILLCELL_X32 FILLER_21_210 ();
 FILLCELL_X8 FILLER_21_242 ();
 FILLCELL_X4 FILLER_21_250 ();
 FILLCELL_X1 FILLER_21_254 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X4 FILLER_22_97 ();
 FILLCELL_X2 FILLER_22_122 ();
 FILLCELL_X2 FILLER_22_133 ();
 FILLCELL_X2 FILLER_22_144 ();
 FILLCELL_X32 FILLER_22_150 ();
 FILLCELL_X32 FILLER_22_182 ();
 FILLCELL_X32 FILLER_22_214 ();
 FILLCELL_X8 FILLER_22_246 ();
 FILLCELL_X1 FILLER_22_254 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X32 FILLER_23_143 ();
 FILLCELL_X32 FILLER_23_175 ();
 FILLCELL_X32 FILLER_23_207 ();
 FILLCELL_X16 FILLER_23_239 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X16 FILLER_24_225 ();
 FILLCELL_X8 FILLER_24_241 ();
 FILLCELL_X4 FILLER_24_249 ();
 FILLCELL_X2 FILLER_24_253 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_97 ();
 FILLCELL_X1 FILLER_25_99 ();
 FILLCELL_X32 FILLER_25_104 ();
 FILLCELL_X32 FILLER_25_136 ();
 FILLCELL_X32 FILLER_25_168 ();
 FILLCELL_X32 FILLER_25_200 ();
 FILLCELL_X16 FILLER_25_232 ();
 FILLCELL_X4 FILLER_25_248 ();
 FILLCELL_X2 FILLER_25_252 ();
 FILLCELL_X1 FILLER_25_254 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X16 FILLER_26_225 ();
 FILLCELL_X8 FILLER_26_241 ();
 FILLCELL_X4 FILLER_26_249 ();
 FILLCELL_X2 FILLER_26_253 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X16 FILLER_27_225 ();
 FILLCELL_X8 FILLER_27_241 ();
 FILLCELL_X4 FILLER_27_249 ();
 FILLCELL_X2 FILLER_27_253 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X16 FILLER_28_225 ();
 FILLCELL_X8 FILLER_28_241 ();
 FILLCELL_X4 FILLER_28_249 ();
 FILLCELL_X2 FILLER_28_253 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X16 FILLER_29_225 ();
 FILLCELL_X8 FILLER_29_241 ();
 FILLCELL_X4 FILLER_29_249 ();
 FILLCELL_X2 FILLER_29_253 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X16 FILLER_30_225 ();
 FILLCELL_X8 FILLER_30_241 ();
 FILLCELL_X4 FILLER_30_249 ();
 FILLCELL_X2 FILLER_30_253 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X16 FILLER_31_225 ();
 FILLCELL_X8 FILLER_31_241 ();
 FILLCELL_X4 FILLER_31_249 ();
 FILLCELL_X2 FILLER_31_253 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X4 FILLER_32_129 ();
 FILLCELL_X2 FILLER_32_133 ();
 FILLCELL_X1 FILLER_32_135 ();
 FILLCELL_X32 FILLER_32_139 ();
 FILLCELL_X32 FILLER_32_171 ();
 FILLCELL_X32 FILLER_32_203 ();
 FILLCELL_X16 FILLER_32_235 ();
 FILLCELL_X4 FILLER_32_251 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_97 ();
 FILLCELL_X4 FILLER_33_113 ();
 FILLCELL_X2 FILLER_33_117 ();
 FILLCELL_X4 FILLER_33_122 ();
 FILLCELL_X2 FILLER_33_126 ();
 FILLCELL_X1 FILLER_33_128 ();
 FILLCELL_X8 FILLER_33_135 ();
 FILLCELL_X2 FILLER_33_143 ();
 FILLCELL_X16 FILLER_33_148 ();
 FILLCELL_X4 FILLER_33_164 ();
 FILLCELL_X2 FILLER_33_168 ();
 FILLCELL_X1 FILLER_33_170 ();
 FILLCELL_X32 FILLER_33_174 ();
 FILLCELL_X32 FILLER_33_206 ();
 FILLCELL_X16 FILLER_33_238 ();
 FILLCELL_X1 FILLER_33_254 ();
endmodule
