module jtag_controller (clk,
    dr_shift_en,
    rst_n,
    tck,
    tdi,
    tdo,
    tms,
    trst_n,
    update_dr,
    dr_in,
    dr_out,
    instruction);
 input clk;
 output dr_shift_en;
 input rst_n;
 input tck;
 input tdi;
 output tdo;
 input tms;
 input trst_n;
 output update_dr;
 input [31:0] dr_in;
 output [31:0] dr_out;
 output [4:0] instruction;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire \dr_shift_reg[0] ;
 wire \dr_shift_reg[10] ;
 wire \dr_shift_reg[11] ;
 wire \dr_shift_reg[12] ;
 wire \dr_shift_reg[13] ;
 wire \dr_shift_reg[14] ;
 wire \dr_shift_reg[15] ;
 wire \dr_shift_reg[16] ;
 wire \dr_shift_reg[17] ;
 wire \dr_shift_reg[18] ;
 wire \dr_shift_reg[19] ;
 wire \dr_shift_reg[1] ;
 wire \dr_shift_reg[20] ;
 wire \dr_shift_reg[21] ;
 wire \dr_shift_reg[22] ;
 wire \dr_shift_reg[23] ;
 wire \dr_shift_reg[24] ;
 wire \dr_shift_reg[25] ;
 wire \dr_shift_reg[26] ;
 wire \dr_shift_reg[27] ;
 wire \dr_shift_reg[28] ;
 wire \dr_shift_reg[29] ;
 wire \dr_shift_reg[2] ;
 wire \dr_shift_reg[30] ;
 wire \dr_shift_reg[31] ;
 wire \dr_shift_reg[3] ;
 wire \dr_shift_reg[4] ;
 wire \dr_shift_reg[5] ;
 wire \dr_shift_reg[6] ;
 wire \dr_shift_reg[7] ;
 wire \dr_shift_reg[8] ;
 wire \dr_shift_reg[9] ;
 wire \ir_shift_reg[0] ;
 wire \ir_shift_reg[1] ;
 wire \ir_shift_reg[2] ;
 wire \ir_shift_reg[3] ;
 wire \ir_shift_reg[4] ;
 wire \next_tap_state[0] ;
 wire \next_tap_state[1] ;
 wire \next_tap_state[2] ;
 wire \next_tap_state[3] ;
 wire \tap_state[0] ;
 wire \tap_state[1] ;
 wire \tap_state[2] ;
 wire \tap_state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _159_ (.I(\tap_state[3] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _160_ (.A1(\tap_state[1] ),
    .A2(\tap_state[0] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _161_ (.A1(_075_),
    .A2(\tap_state[2] ),
    .A3(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _162_ (.I(_077_),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _163_ (.A1(\dr_shift_reg[0] ),
    .A2(net69),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _164_ (.I(\tap_state[1] ),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _165_ (.I(\tap_state[0] ),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _166_ (.I(\tap_state[2] ),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _167_ (.A1(\tap_state[3] ),
    .A2(_081_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _168_ (.A1(_079_),
    .A2(_080_),
    .A3(\ir_shift_reg[0] ),
    .A4(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _169_ (.A1(_078_),
    .A2(_083_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _170_ (.A1(_076_),
    .A2(_082_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _171_ (.I(_084_),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _172_ (.I0(net52),
    .I1(\dr_shift_reg[23] ),
    .S(net76),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _173_ (.I0(net53),
    .I1(\dr_shift_reg[24] ),
    .S(net76),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _174_ (.I0(net54),
    .I1(\dr_shift_reg[25] ),
    .S(net76),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _175_ (.I0(net55),
    .I1(\dr_shift_reg[26] ),
    .S(net76),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _176_ (.I0(net56),
    .I1(\dr_shift_reg[27] ),
    .S(net76),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _177_ (.I0(net57),
    .I1(\dr_shift_reg[28] ),
    .S(net76),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _178_ (.I0(net58),
    .I1(\dr_shift_reg[29] ),
    .S(net76),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _179_ (.I0(net59),
    .I1(\dr_shift_reg[2] ),
    .S(net76),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _180_ (.I0(net60),
    .I1(\dr_shift_reg[30] ),
    .S(net76),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _181_ (.I(_084_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _182_ (.I0(net61),
    .I1(\dr_shift_reg[31] ),
    .S(_085_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _183_ (.I0(net62),
    .I1(\dr_shift_reg[3] ),
    .S(_085_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _184_ (.I0(net63),
    .I1(\dr_shift_reg[4] ),
    .S(_085_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _185_ (.I0(net64),
    .I1(\dr_shift_reg[5] ),
    .S(_085_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _186_ (.I0(net65),
    .I1(\dr_shift_reg[6] ),
    .S(_085_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _187_ (.I0(net66),
    .I1(\dr_shift_reg[7] ),
    .S(_085_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _188_ (.I0(net67),
    .I1(\dr_shift_reg[8] ),
    .S(_085_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _189_ (.I0(net68),
    .I1(\dr_shift_reg[9] ),
    .S(_085_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _190_ (.I(\dr_shift_reg[0] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _191_ (.A1(\tap_state[3] ),
    .A2(\tap_state[2] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _192_ (.A1(\tap_state[1] ),
    .A2(\tap_state[0] ),
    .A3(_087_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _193_ (.A1(_077_),
    .A2(_088_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _194_ (.I(_089_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _195_ (.I(_088_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _196_ (.I(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _197_ (.A1(\dr_shift_reg[1] ),
    .A2(net69),
    .B1(_092_),
    .B2(net1),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _198_ (.A1(_086_),
    .A2(_090_),
    .B(_093_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _199_ (.I(\dr_shift_reg[10] ),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _200_ (.A1(\dr_shift_reg[11] ),
    .A2(net69),
    .B1(_092_),
    .B2(net2),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _201_ (.A1(_094_),
    .A2(_090_),
    .B(_095_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _202_ (.I(\dr_shift_reg[11] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _203_ (.A1(\dr_shift_reg[12] ),
    .A2(net69),
    .B1(_092_),
    .B2(net3),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _204_ (.A1(_096_),
    .A2(_090_),
    .B(_097_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _205_ (.I0(\dr_shift_reg[13] ),
    .I1(net4),
    .S(_091_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _206_ (.I0(\dr_shift_reg[12] ),
    .I1(_098_),
    .S(_090_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _207_ (.I0(\dr_shift_reg[13] ),
    .I1(\dr_shift_reg[14] ),
    .S(net69),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _208_ (.I0(_099_),
    .I1(net5),
    .S(_092_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(\dr_shift_reg[15] ),
    .I1(net6),
    .S(_091_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _210_ (.I0(\dr_shift_reg[14] ),
    .I1(_100_),
    .S(_090_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(\dr_shift_reg[16] ),
    .I1(net7),
    .S(_091_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(\dr_shift_reg[15] ),
    .I1(_101_),
    .S(_090_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _213_ (.I0(\dr_shift_reg[16] ),
    .I1(\dr_shift_reg[17] ),
    .S(net69),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(_102_),
    .I1(net8),
    .S(_092_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(\dr_shift_reg[18] ),
    .I1(net9),
    .S(_091_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(\dr_shift_reg[17] ),
    .I1(_103_),
    .S(_090_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _217_ (.I(\dr_shift_reg[18] ),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _218_ (.A1(\dr_shift_reg[19] ),
    .A2(net69),
    .B1(_092_),
    .B2(net10),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _219_ (.A1(_104_),
    .A2(_090_),
    .B(_105_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _220_ (.I0(\dr_shift_reg[20] ),
    .I1(net11),
    .S(_091_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(\dr_shift_reg[19] ),
    .I1(_106_),
    .S(_090_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _222_ (.I0(\dr_shift_reg[1] ),
    .I1(\dr_shift_reg[2] ),
    .S(net69),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(_107_),
    .I1(net12),
    .S(_092_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(\dr_shift_reg[21] ),
    .I1(net13),
    .S(_091_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _225_ (.I0(\dr_shift_reg[20] ),
    .I1(_108_),
    .S(_090_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(\dr_shift_reg[22] ),
    .I1(net14),
    .S(_091_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _227_ (.I(_089_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _228_ (.I0(\dr_shift_reg[21] ),
    .I1(_109_),
    .S(_110_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _229_ (.I0(\dr_shift_reg[23] ),
    .I1(net15),
    .S(_091_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _230_ (.I0(\dr_shift_reg[22] ),
    .I1(_111_),
    .S(_110_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _231_ (.I(_088_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _232_ (.I0(\dr_shift_reg[24] ),
    .I1(net16),
    .S(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(\dr_shift_reg[23] ),
    .I1(_113_),
    .S(_110_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _234_ (.I0(\dr_shift_reg[24] ),
    .I1(\dr_shift_reg[25] ),
    .S(net69),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _235_ (.I0(_114_),
    .I1(net17),
    .S(_092_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _236_ (.I0(\dr_shift_reg[26] ),
    .I1(net18),
    .S(_112_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _237_ (.I0(\dr_shift_reg[25] ),
    .I1(_115_),
    .S(_110_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(\dr_shift_reg[26] ),
    .I1(\dr_shift_reg[27] ),
    .S(_077_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _239_ (.I0(_116_),
    .I1(net19),
    .S(_092_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(\dr_shift_reg[28] ),
    .I1(net20),
    .S(_112_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _241_ (.I0(\dr_shift_reg[27] ),
    .I1(_117_),
    .S(_110_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _242_ (.I0(\dr_shift_reg[29] ),
    .I1(net21),
    .S(_112_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _243_ (.I0(\dr_shift_reg[28] ),
    .I1(_118_),
    .S(_110_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(\dr_shift_reg[30] ),
    .I1(net22),
    .S(_112_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _245_ (.I0(\dr_shift_reg[29] ),
    .I1(_119_),
    .S(_110_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _246_ (.I0(\dr_shift_reg[3] ),
    .I1(net23),
    .S(_112_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _247_ (.I0(\dr_shift_reg[2] ),
    .I1(_120_),
    .S(_110_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _248_ (.I0(\dr_shift_reg[31] ),
    .I1(net24),
    .S(_112_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _249_ (.I0(\dr_shift_reg[30] ),
    .I1(_121_),
    .S(_110_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _250_ (.I0(net34),
    .I1(net25),
    .S(_112_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _251_ (.I0(\dr_shift_reg[31] ),
    .I1(_122_),
    .S(_110_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _252_ (.I0(\dr_shift_reg[3] ),
    .I1(\dr_shift_reg[4] ),
    .S(_077_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _253_ (.I0(_123_),
    .I1(net26),
    .S(_092_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _254_ (.I0(\dr_shift_reg[4] ),
    .I1(\dr_shift_reg[5] ),
    .S(_077_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _255_ (.I0(_124_),
    .I1(net27),
    .S(_091_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _256_ (.I0(\dr_shift_reg[6] ),
    .I1(net28),
    .S(_112_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _257_ (.I0(\dr_shift_reg[5] ),
    .I1(_125_),
    .S(_089_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _258_ (.I0(\dr_shift_reg[7] ),
    .I1(net29),
    .S(_112_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _259_ (.I0(\dr_shift_reg[6] ),
    .I1(_126_),
    .S(_089_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _260_ (.I0(\dr_shift_reg[8] ),
    .I1(net30),
    .S(_088_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _261_ (.I0(\dr_shift_reg[7] ),
    .I1(_127_),
    .S(_089_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _262_ (.I0(\dr_shift_reg[9] ),
    .I1(net31),
    .S(_088_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _263_ (.I0(\dr_shift_reg[8] ),
    .I1(_128_),
    .S(_089_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _264_ (.I0(\dr_shift_reg[10] ),
    .I1(net32),
    .S(_088_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _265_ (.I0(\dr_shift_reg[9] ),
    .I1(_129_),
    .S(_089_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _266_ (.I(_080_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _267_ (.A1(_130_),
    .A2(\ir_shift_reg[1] ),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _268_ (.A1(_079_),
    .A2(_082_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _269_ (.I0(\ir_shift_reg[0] ),
    .I1(_131_),
    .S(_132_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _270_ (.A1(_130_),
    .A2(\ir_shift_reg[2] ),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _271_ (.I0(\ir_shift_reg[1] ),
    .I1(_133_),
    .S(_132_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _272_ (.A1(_130_),
    .A2(\ir_shift_reg[3] ),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _273_ (.I0(\ir_shift_reg[2] ),
    .I1(_134_),
    .S(_132_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _274_ (.A1(_130_),
    .A2(\ir_shift_reg[4] ),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _275_ (.I0(\ir_shift_reg[3] ),
    .I1(_135_),
    .S(_132_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _276_ (.A1(_080_),
    .A2(net34),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _277_ (.I0(\ir_shift_reg[4] ),
    .I1(_136_),
    .S(_132_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _278_ (.I0(net37),
    .I1(\dr_shift_reg[0] ),
    .S(_085_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _279_ (.I0(net38),
    .I1(\dr_shift_reg[10] ),
    .S(_085_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _280_ (.I(_084_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _281_ (.I0(net39),
    .I1(\dr_shift_reg[11] ),
    .S(_137_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _282_ (.I0(net40),
    .I1(\dr_shift_reg[12] ),
    .S(_137_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _283_ (.I0(net41),
    .I1(\dr_shift_reg[13] ),
    .S(_137_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _284_ (.I0(net42),
    .I1(\dr_shift_reg[14] ),
    .S(_137_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _285_ (.I0(net43),
    .I1(\dr_shift_reg[15] ),
    .S(_137_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _286_ (.I0(net44),
    .I1(\dr_shift_reg[16] ),
    .S(_137_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _287_ (.I0(net45),
    .I1(\dr_shift_reg[17] ),
    .S(_137_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _288_ (.I0(net46),
    .I1(\dr_shift_reg[18] ),
    .S(_137_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _289_ (.I0(net47),
    .I1(\dr_shift_reg[19] ),
    .S(_137_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _290_ (.I0(net48),
    .I1(\dr_shift_reg[1] ),
    .S(_137_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _291_ (.I0(net49),
    .I1(\dr_shift_reg[20] ),
    .S(_084_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _292_ (.I0(net50),
    .I1(\dr_shift_reg[21] ),
    .S(_084_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _293_ (.I0(net51),
    .I1(\dr_shift_reg[22] ),
    .S(_084_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _294_ (.A1(\tap_state[1] ),
    .A2(_080_),
    .A3(\tap_state[3] ),
    .A4(\tap_state[2] ),
    .Z(_138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _295_ (.I0(net70),
    .I1(\ir_shift_reg[0] ),
    .S(_138_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _296_ (.I0(net71),
    .I1(\ir_shift_reg[1] ),
    .S(_138_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _297_ (.I0(net72),
    .I1(\ir_shift_reg[2] ),
    .S(_138_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _298_ (.I0(net73),
    .I1(\ir_shift_reg[3] ),
    .S(_138_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _299_ (.I0(net74),
    .I1(\ir_shift_reg[4] ),
    .S(_138_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _300_ (.I(net35),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _301_ (.A1(_079_),
    .A2(_139_),
    .B(\tap_state[2] ),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _302_ (.A1(_081_),
    .A2(net35),
    .B1(_140_),
    .B2(_130_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _303_ (.A1(_080_),
    .A2(\tap_state[3] ),
    .B(net35),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _304_ (.A1(_080_),
    .A2(_081_),
    .B(net35),
    .C(\tap_state[3] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _305_ (.A1(_079_),
    .A2(\tap_state[2] ),
    .A3(_142_),
    .B(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _306_ (.A1(_075_),
    .A2(_141_),
    .B(_144_),
    .ZN(\next_tap_state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _307_ (.A1(_079_),
    .A2(\tap_state[3] ),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _308_ (.A1(\tap_state[2] ),
    .A2(net35),
    .Z(_146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _309_ (.A1(_139_),
    .A2(_082_),
    .B1(_145_),
    .B2(_146_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _310_ (.A1(\tap_state[3] ),
    .A2(net35),
    .B(_079_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _311_ (.A1(_079_),
    .A2(_081_),
    .A3(net35),
    .Z(_149_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _312_ (.A1(_080_),
    .A2(_148_),
    .A3(_149_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _313_ (.A1(_075_),
    .A2(_081_),
    .A3(_139_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _314_ (.A1(_130_),
    .A2(_147_),
    .B(_150_),
    .C(_151_),
    .ZN(\next_tap_state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _315_ (.A1(_130_),
    .A2(_081_),
    .A3(_139_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _316_ (.A1(_075_),
    .A2(net35),
    .B(_152_),
    .C(_079_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _317_ (.A1(_080_),
    .A2(_075_),
    .A3(net35),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _318_ (.A1(_079_),
    .A2(_081_),
    .A3(_154_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _319_ (.A1(_130_),
    .A2(_087_),
    .B1(_153_),
    .B2(_155_),
    .ZN(\next_tap_state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _320_ (.A1(_080_),
    .A2(_139_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _321_ (.A1(_130_),
    .A2(\tap_state[3] ),
    .B1(_156_),
    .B2(_079_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _322_ (.A1(_080_),
    .A2(_081_),
    .B(net35),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _323_ (.A1(_081_),
    .A2(_157_),
    .B1(_158_),
    .B2(_075_),
    .C(_138_),
    .ZN(\next_tap_state[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[0]$_DFFE_NN0P_  (.D(_060_),
    .RN(net36),
    .CLKN(net33),
    .Q(net37));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[10]$_DFFE_NN0P_  (.D(_061_),
    .RN(net36),
    .CLKN(net33),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[11]$_DFFE_NN0P_  (.D(_062_),
    .RN(net36),
    .CLKN(net33),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[12]$_DFFE_NN0P_  (.D(_063_),
    .RN(net36),
    .CLKN(net33),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[13]$_DFFE_NN0P_  (.D(_064_),
    .RN(net36),
    .CLKN(net33),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[14]$_DFFE_NN0P_  (.D(_065_),
    .RN(net36),
    .CLKN(net33),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[15]$_DFFE_NN0P_  (.D(_066_),
    .RN(net36),
    .CLKN(net33),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[16]$_DFFE_NN0P_  (.D(_067_),
    .RN(net36),
    .CLKN(net33),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[17]$_DFFE_NN0P_  (.D(_068_),
    .RN(net36),
    .CLKN(net33),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[18]$_DFFE_NN0P_  (.D(_069_),
    .RN(net36),
    .CLKN(net33),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[19]$_DFFE_NN0P_  (.D(_070_),
    .RN(net36),
    .CLKN(net33),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[1]$_DFFE_NN0P_  (.D(_071_),
    .RN(net36),
    .CLKN(net33),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[20]$_DFFE_NN0P_  (.D(_072_),
    .RN(net36),
    .CLKN(net33),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[21]$_DFFE_NN0P_  (.D(_073_),
    .RN(net36),
    .CLKN(net33),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[22]$_DFFE_NN0P_  (.D(_074_),
    .RN(net36),
    .CLKN(net33),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[23]$_DFFE_NN0P_  (.D(_001_),
    .RN(net36),
    .CLKN(net33),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[24]$_DFFE_NN0P_  (.D(_002_),
    .RN(net36),
    .CLKN(net33),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[25]$_DFFE_NN0P_  (.D(_003_),
    .RN(net36),
    .CLKN(net33),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[26]$_DFFE_NN0P_  (.D(_004_),
    .RN(net36),
    .CLKN(net33),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[27]$_DFFE_NN0P_  (.D(_005_),
    .RN(net36),
    .CLKN(net33),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[28]$_DFFE_NN0P_  (.D(_006_),
    .RN(net36),
    .CLKN(net33),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[29]$_DFFE_NN0P_  (.D(_007_),
    .RN(net36),
    .CLKN(net33),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[2]$_DFFE_NN0P_  (.D(_008_),
    .RN(net36),
    .CLKN(net33),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[30]$_DFFE_NN0P_  (.D(_009_),
    .RN(net36),
    .CLKN(net33),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[31]$_DFFE_NN0P_  (.D(_010_),
    .RN(net36),
    .CLKN(net33),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[3]$_DFFE_NN0P_  (.D(_011_),
    .RN(net36),
    .CLKN(net33),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[4]$_DFFE_NN0P_  (.D(_012_),
    .RN(net36),
    .CLKN(net33),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[5]$_DFFE_NN0P_  (.D(_013_),
    .RN(net36),
    .CLKN(net33),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[6]$_DFFE_NN0P_  (.D(_014_),
    .RN(net36),
    .CLKN(net33),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[7]$_DFFE_NN0P_  (.D(_015_),
    .RN(net36),
    .CLKN(net33),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[8]$_DFFE_NN0P_  (.D(_016_),
    .RN(net36),
    .CLKN(net33),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \dr_reg[9]$_DFFE_NN0P_  (.D(_017_),
    .RN(net36),
    .CLKN(net33),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[0]$_DFFE_PN0P_  (.D(_018_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[10]$_DFFE_PN0P_  (.D(_019_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[11]$_DFFE_PN0P_  (.D(_020_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[12]$_DFFE_PN0P_  (.D(_021_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[13]$_DFFE_PN0P_  (.D(_022_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[14]$_DFFE_PN0P_  (.D(_023_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[15]$_DFFE_PN0P_  (.D(_024_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[16]$_DFFE_PN0P_  (.D(_025_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[17]$_DFFE_PN0P_  (.D(_026_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[18]$_DFFE_PN0P_  (.D(_027_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[19]$_DFFE_PN0P_  (.D(_028_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[1]$_DFFE_PN0P_  (.D(_029_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[20]$_DFFE_PN0P_  (.D(_030_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[21]$_DFFE_PN0P_  (.D(_031_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[22]$_DFFE_PN0P_  (.D(_032_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[23]$_DFFE_PN0P_  (.D(_033_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[24]$_DFFE_PN0P_  (.D(_034_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[25]$_DFFE_PN0P_  (.D(_035_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[26]$_DFFE_PN0P_  (.D(_036_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[27]$_DFFE_PN0P_  (.D(_037_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[28]$_DFFE_PN0P_  (.D(_038_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[29]$_DFFE_PN0P_  (.D(_039_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[2]$_DFFE_PN0P_  (.D(_040_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[30]$_DFFE_PN0P_  (.D(_041_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[31]$_DFFE_PN0P_  (.D(_042_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[3]$_DFFE_PN0P_  (.D(_043_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[4]$_DFFE_PN0P_  (.D(_044_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[5]$_DFFE_PN0P_  (.D(_045_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[6]$_DFFE_PN0P_  (.D(_046_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[7]$_DFFE_PN0P_  (.D(_047_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[8]$_DFFE_PN0P_  (.D(_048_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dr_shift_reg[9]$_DFFE_PN0P_  (.D(_049_),
    .RN(net36),
    .CLK(net33),
    .Q(\dr_shift_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 \ir_reg[0]$_DFFE_NN1N_  (.D(_050_),
    .SETN(net36),
    .CLKN(net33),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \ir_reg[1]$_DFFE_NN0N_  (.D(_051_),
    .RN(net36),
    .CLKN(net33),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \ir_reg[2]$_DFFE_NN0N_  (.D(_052_),
    .RN(net36),
    .CLKN(net33),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \ir_reg[3]$_DFFE_NN0N_  (.D(_053_),
    .RN(net36),
    .CLKN(net33),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \ir_reg[4]$_DFFE_NN0N_  (.D(_054_),
    .RN(net36),
    .CLKN(net33),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \ir_shift_reg[0]$_DFFE_PN1P_  (.D(_055_),
    .SETN(net36),
    .CLK(net33),
    .Q(\ir_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ir_shift_reg[1]$_DFFE_PN0P_  (.D(_056_),
    .RN(net36),
    .CLK(net33),
    .Q(\ir_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ir_shift_reg[2]$_DFFE_PN0P_  (.D(_057_),
    .RN(net36),
    .CLK(net33),
    .Q(\ir_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ir_shift_reg[3]$_DFFE_PN0P_  (.D(_058_),
    .RN(net36),
    .CLK(net33),
    .Q(\ir_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ir_shift_reg[4]$_DFFE_PN0P_  (.D(_059_),
    .RN(net36),
    .CLK(net33),
    .Q(\ir_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tap_state[0]$_DFF_PN0_  (.D(\next_tap_state[0] ),
    .RN(net36),
    .CLK(net33),
    .Q(\tap_state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tap_state[1]$_DFF_PN0_  (.D(\next_tap_state[1] ),
    .RN(net36),
    .CLK(net33),
    .Q(\tap_state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tap_state[2]$_DFF_PN0_  (.D(\next_tap_state[2] ),
    .RN(net36),
    .CLK(net33),
    .Q(\tap_state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \tap_state[3]$_DFF_PN0_  (.D(\next_tap_state[3] ),
    .RN(net36),
    .CLK(net33),
    .Q(\tap_state[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 \tdo_mux$_DFF_NN0_  (.D(_000_),
    .RN(net36),
    .CLKN(net33),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_77 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_78 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_79 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_80 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_90 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(dr_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(dr_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(dr_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(dr_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(dr_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(dr_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(dr_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(dr_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(dr_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(dr_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(dr_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(dr_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(dr_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(dr_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(dr_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(dr_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(dr_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(dr_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(dr_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(dr_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(dr_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(dr_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(dr_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(dr_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(dr_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(dr_in[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(dr_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(dr_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(dr_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(dr_in[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(dr_in[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(dr_in[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 input33 (.I(tck),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(tdi),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input35 (.I(tms),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input36 (.I(trst_n),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net37),
    .Z(dr_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net38),
    .Z(dr_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net39),
    .Z(dr_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net40),
    .Z(dr_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net41),
    .Z(dr_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net42),
    .Z(dr_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net43),
    .Z(dr_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net44),
    .Z(dr_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net45),
    .Z(dr_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net46),
    .Z(dr_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net47),
    .Z(dr_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net48),
    .Z(dr_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net49),
    .Z(dr_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net50),
    .Z(dr_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net51),
    .Z(dr_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net52),
    .Z(dr_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net53),
    .Z(dr_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net54),
    .Z(dr_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net55),
    .Z(dr_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net56),
    .Z(dr_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net57),
    .Z(dr_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net58),
    .Z(dr_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net59),
    .Z(dr_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net60),
    .Z(dr_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net61),
    .Z(dr_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net62),
    .Z(dr_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net63),
    .Z(dr_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net64),
    .Z(dr_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net65),
    .Z(dr_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(dr_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(dr_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(dr_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(dr_shift_en));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(instruction[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(instruction[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(instruction[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(instruction[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(instruction[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(tdo));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(update_dr));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_333 ();
endmodule
