module fair_priority_arbiter (clk,
    rst_n,
    valid,
    grant,
    grant_idx,
    priorities,
    request);
 input clk;
 input rst_n;
 output valid;
 output [3:0] grant;
 output [1:0] grant_idx;
 input [7:0] priorities;
 input [3:0] request;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire net53;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;

 CLKBUF_X3 _184_ (.A(_152_),
    .Z(_100_));
 CLKBUF_X3 _185_ (.A(_164_),
    .Z(_101_));
 BUF_X1 rebuffer37 (.A(_016_),
    .Z(net53));
 AOI222_X2 _187_ (.A1(net5),
    .A2(_100_),
    .B1(_101_),
    .B2(net3),
    .C1(_160_),
    .C2(net7),
    .ZN(_103_));
 INV_X1 _188_ (.A(_103_),
    .ZN(_104_));
 MUX2_X1 _189_ (.A(_104_),
    .B(net1),
    .S(_158_),
    .Z(_105_));
 INV_X1 _190_ (.A(_105_),
    .ZN(_147_));
 AOI222_X2 _191_ (.A1(net6),
    .A2(_100_),
    .B1(_101_),
    .B2(net4),
    .C1(_160_),
    .C2(net8),
    .ZN(_106_));
 INV_X1 _192_ (.A(net2),
    .ZN(_107_));
 MUX2_X1 _193_ (.A(_106_),
    .B(_107_),
    .S(_158_),
    .Z(_108_));
 INV_X1 _194_ (.A(_108_),
    .ZN(_143_));
 CLKBUF_X3 _195_ (.A(_156_),
    .Z(_109_));
 AOI222_X2 _196_ (.A1(net7),
    .A2(_100_),
    .B1(_109_),
    .B2(net3),
    .C1(_101_),
    .C2(net5),
    .ZN(_110_));
 INV_X1 _197_ (.A(_110_),
    .ZN(_111_));
 MUX2_X1 _198_ (.A(_111_),
    .B(net1),
    .S(_162_),
    .Z(_112_));
 INV_X1 _199_ (.A(_112_),
    .ZN(_173_));
 AOI222_X2 _200_ (.A1(net8),
    .A2(_100_),
    .B1(_109_),
    .B2(net4),
    .C1(_101_),
    .C2(net6),
    .ZN(_113_));
 MUX2_X1 _201_ (.A(_113_),
    .B(_107_),
    .S(_162_),
    .Z(_114_));
 INV_X1 _202_ (.A(_114_),
    .ZN(_169_));
 AOI222_X2 _203_ (.A1(net5),
    .A2(_109_),
    .B1(_160_),
    .B2(net3),
    .C1(_101_),
    .C2(net7),
    .ZN(_115_));
 INV_X1 _204_ (.A(net1),
    .ZN(_116_));
 MUX2_X1 _205_ (.A(_115_),
    .B(_116_),
    .S(_154_),
    .Z(_180_));
 BUF_X4 _206_ (.A(_166_),
    .Z(_117_));
 BUF_X4 _207_ (.A(request[0]),
    .Z(_118_));
 BUF_X4 _208_ (.A(request[2]),
    .Z(_119_));
 MUX2_X1 _209_ (.A(_118_),
    .B(_119_),
    .S(net18),
    .Z(_120_));
 AND3_X1 _210_ (.A1(_117_),
    .A2(net2),
    .A3(_120_),
    .ZN(_121_));
 CLKBUF_X3 _211_ (.A(request[1]),
    .Z(_122_));
 CLKBUF_X3 _212_ (.A(request[3]),
    .Z(_123_));
 BUF_X4 _213_ (.A(_153_),
    .Z(_124_));
 MUX2_X2 _214_ (.A(_122_),
    .B(_123_),
    .S(_124_),
    .Z(_125_));
 BUF_X4 _215_ (.A(net14),
    .Z(_126_));
 MUX2_X1 _216_ (.A(_125_),
    .B(_120_),
    .S(_126_),
    .Z(_127_));
 AOI222_X2 _217_ (.A1(net8),
    .A2(_109_),
    .B1(_160_),
    .B2(net6),
    .C1(net4),
    .C2(_100_),
    .ZN(_128_));
 NOR2_X1 _218_ (.A1(_117_),
    .A2(_128_),
    .ZN(_129_));
 AOI21_X2 _219_ (.A(_121_),
    .B1(_127_),
    .B2(_129_),
    .ZN(_142_));
 NAND3_X1 _220_ (.A1(_117_),
    .A2(net1),
    .A3(net37),
    .ZN(_130_));
 AOI222_X2 _221_ (.A1(net7),
    .A2(_109_),
    .B1(_160_),
    .B2(net5),
    .C1(net3),
    .C2(_100_),
    .ZN(_131_));
 INV_X1 _222_ (.A(_131_),
    .ZN(_132_));
 NAND2_X1 _223_ (.A1(_127_),
    .A2(_132_),
    .ZN(_133_));
 OAI21_X1 _224_ (.A(_130_),
    .B1(_133_),
    .B2(_117_),
    .ZN(_146_));
 OR2_X1 _225_ (.A1(_117_),
    .A2(_126_),
    .ZN(_134_));
 BUF_X8 _226_ (.A(_134_),
    .Z(_135_));
 MUX2_X1 _227_ (.A(_119_),
    .B(_118_),
    .S(net19),
    .Z(_136_));
 NOR2_X1 _228_ (.A1(_135_),
    .A2(_136_),
    .ZN(_007_));
 INV_X1 _229_ (.A(_007_),
    .ZN(_008_));
 NOR2_X4 _230_ (.A1(_117_),
    .A2(_126_),
    .ZN(_009_));
 CLKBUF_X3 _231_ (.A(_009_),
    .Z(_010_));
 OAI21_X1 _232_ (.A(_008_),
    .B1(_010_),
    .B2(net34),
    .ZN(_011_));
 NOR2_X1 _233_ (.A1(net38),
    .A2(_009_),
    .ZN(_012_));
 NAND2_X2 _234_ (.A1(net20),
    .A2(_149_),
    .ZN(_013_));
 INV_X1 _235_ (.A(_144_),
    .ZN(_014_));
 INV_X1 _236_ (.A(_145_),
    .ZN(_015_));
 OAI21_X4 _237_ (.A(_014_),
    .B1(_015_),
    .B2(_148_),
    .ZN(_016_));
 AOI21_X2 _238_ (.A(_012_),
    .B1(_013_),
    .B2(_016_),
    .ZN(_017_));
 AOI21_X2 _239_ (.A(_011_),
    .B1(_017_),
    .B2(net35),
    .ZN(_018_));
 MUX2_X1 _240_ (.A(_142_),
    .B(_108_),
    .S(_018_),
    .Z(_168_));
 MUX2_X1 _241_ (.A(_146_),
    .B(_105_),
    .S(_018_),
    .Z(_172_));
 MUX2_X1 _242_ (.A(_123_),
    .B(_122_),
    .S(net23),
    .Z(_019_));
 OR2_X1 _243_ (.A1(_135_),
    .A2(_019_),
    .ZN(_020_));
 OAI21_X2 _244_ (.A(_020_),
    .B1(_136_),
    .B2(_010_),
    .ZN(_021_));
 INV_X1 _245_ (.A(_174_),
    .ZN(_022_));
 AOI21_X2 _246_ (.A(_170_),
    .B1(_022_),
    .B2(_171_),
    .ZN(_023_));
 AOI21_X4 _247_ (.A(_023_),
    .B1(_175_),
    .B2(net17),
    .ZN(_024_));
 NOR3_X2 _248_ (.A1(_117_),
    .A2(_126_),
    .A3(_123_),
    .ZN(_025_));
 NOR2_X2 _249_ (.A1(_122_),
    .A2(net24),
    .ZN(_026_));
 AOI22_X4 _250_ (.A1(net25),
    .A2(_025_),
    .B1(_026_),
    .B2(_135_),
    .ZN(_027_));
 NOR2_X4 _251_ (.A1(_118_),
    .A2(_027_),
    .ZN(_028_));
 INV_X1 _252_ (.A(_123_),
    .ZN(_029_));
 NAND3_X2 _253_ (.A1(_029_),
    .A2(net26),
    .A3(_135_),
    .ZN(_030_));
 NAND2_X1 _254_ (.A1(_009_),
    .A2(_026_),
    .ZN(_031_));
 AOI21_X4 _255_ (.A(_119_),
    .B1(_030_),
    .B2(_031_),
    .ZN(_032_));
 NOR3_X4 _256_ (.A1(_024_),
    .A2(_028_),
    .A3(_032_),
    .ZN(_033_));
 NOR2_X4 _257_ (.A1(_033_),
    .A2(_021_),
    .ZN(_034_));
 MUX2_X1 _258_ (.A(_168_),
    .B(_114_),
    .S(_034_),
    .Z(_176_));
 AOI222_X2 _259_ (.A1(net6),
    .A2(_109_),
    .B1(_160_),
    .B2(net4),
    .C1(_101_),
    .C2(net8),
    .ZN(_035_));
 INV_X1 _260_ (.A(_035_),
    .ZN(_036_));
 MUX2_X1 _261_ (.A(_036_),
    .B(net2),
    .S(_154_),
    .Z(_177_));
 MUX2_X1 _262_ (.A(_172_),
    .B(_112_),
    .S(_034_),
    .Z(_181_));
 MUX2_X1 _263_ (.A(_122_),
    .B(_119_),
    .S(_009_),
    .Z(_037_));
 MUX2_X1 _264_ (.A(_118_),
    .B(_123_),
    .S(_135_),
    .Z(_038_));
 INV_X1 _265_ (.A(net26),
    .ZN(_039_));
 MUX2_X1 _266_ (.A(_037_),
    .B(_038_),
    .S(_039_),
    .Z(_040_));
 MUX2_X2 _267_ (.A(_136_),
    .B(_019_),
    .S(_009_),
    .Z(_041_));
 INV_X1 _268_ (.A(_182_),
    .ZN(_042_));
 AOI21_X2 _269_ (.A(_178_),
    .B1(_042_),
    .B2(_179_),
    .ZN(_043_));
 AND2_X2 _270_ (.A1(_179_),
    .A2(_183_),
    .ZN(_044_));
 OAI21_X1 _271_ (.A(_041_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_045_));
 NAND2_X1 _272_ (.A1(_040_),
    .A2(_045_),
    .ZN(_046_));
 NOR2_X2 _273_ (.A1(_043_),
    .A2(_044_),
    .ZN(_047_));
 NOR3_X4 _274_ (.A1(_047_),
    .A2(_032_),
    .A3(_028_),
    .ZN(_048_));
 NOR3_X1 _275_ (.A1(_010_),
    .A2(_046_),
    .A3(_048_),
    .ZN(_049_));
 INV_X1 _276_ (.A(net35),
    .ZN(_050_));
 OR3_X1 _277_ (.A1(_050_),
    .A2(_010_),
    .A3(_017_),
    .ZN(_051_));
 OR3_X2 _278_ (.A1(_024_),
    .A2(_028_),
    .A3(_032_),
    .ZN(_052_));
 AOI21_X1 _279_ (.A(_051_),
    .B1(_052_),
    .B2(_041_),
    .ZN(_053_));
 INV_X1 _280_ (.A(_148_),
    .ZN(_054_));
 AOI21_X2 _281_ (.A(_144_),
    .B1(_054_),
    .B2(net20),
    .ZN(_055_));
 AND2_X1 _282_ (.A1(net21),
    .A2(_149_),
    .ZN(_056_));
 NOR4_X2 _283_ (.A1(_050_),
    .A2(_007_),
    .A3(_055_),
    .A4(_056_),
    .ZN(_057_));
 NOR2_X1 _284_ (.A1(net36),
    .A2(_135_),
    .ZN(_058_));
 OR2_X1 _285_ (.A1(_012_),
    .A2(_058_),
    .ZN(_059_));
 OAI22_X2 _286_ (.A1(_021_),
    .A2(_033_),
    .B1(_057_),
    .B2(_059_),
    .ZN(_060_));
 AND2_X2 _287_ (.A1(_040_),
    .A2(_045_),
    .ZN(_061_));
 OR3_X4 _288_ (.A1(_028_),
    .A2(_032_),
    .A3(_047_),
    .ZN(_062_));
 AOI21_X4 _289_ (.A(_135_),
    .B1(_061_),
    .B2(_062_),
    .ZN(_063_));
 AOI211_X2 _290_ (.A(_049_),
    .B(_053_),
    .C1(_060_),
    .C2(_063_),
    .ZN(_064_));
 NAND3_X1 _291_ (.A1(_122_),
    .A2(net24),
    .A3(_135_),
    .ZN(_065_));
 NAND3_X1 _292_ (.A1(_118_),
    .A2(_039_),
    .A3(_010_),
    .ZN(_066_));
 NAND2_X1 _293_ (.A1(_065_),
    .A2(_066_),
    .ZN(_067_));
 OR2_X1 _294_ (.A1(_118_),
    .A2(_027_),
    .ZN(_068_));
 INV_X1 _295_ (.A(_119_),
    .ZN(_069_));
 NOR3_X1 _296_ (.A1(_123_),
    .A2(_039_),
    .A3(_010_),
    .ZN(_070_));
 AND2_X1 _297_ (.A1(_010_),
    .A2(_026_),
    .ZN(_071_));
 OAI21_X1 _298_ (.A(_069_),
    .B1(_070_),
    .B2(_071_),
    .ZN(_072_));
 AOI21_X1 _299_ (.A(_041_),
    .B1(_068_),
    .B2(_072_),
    .ZN(_073_));
 OAI21_X1 _300_ (.A(_067_),
    .B1(_073_),
    .B2(_047_),
    .ZN(_074_));
 INV_X1 _301_ (.A(_118_),
    .ZN(_075_));
 AOI21_X1 _302_ (.A(_075_),
    .B1(net53),
    .B2(_013_),
    .ZN(_076_));
 NAND3_X1 _303_ (.A1(_122_),
    .A2(_039_),
    .A3(_135_),
    .ZN(_077_));
 AOI21_X1 _304_ (.A(_029_),
    .B1(net53),
    .B2(_013_),
    .ZN(_078_));
 NAND3_X1 _305_ (.A1(_118_),
    .A2(net27),
    .A3(_010_),
    .ZN(_079_));
 OAI22_X2 _306_ (.A1(_076_),
    .A2(_077_),
    .B1(_078_),
    .B2(_079_),
    .ZN(_080_));
 MUX2_X1 _307_ (.A(_119_),
    .B(_123_),
    .S(_009_),
    .Z(_081_));
 NAND2_X1 _308_ (.A1(net28),
    .A2(_081_),
    .ZN(_082_));
 MUX2_X1 _309_ (.A(_118_),
    .B(_122_),
    .S(_009_),
    .Z(_083_));
 OAI21_X1 _310_ (.A(_083_),
    .B1(_056_),
    .B2(_055_),
    .ZN(_084_));
 OAI221_X2 _311_ (.A(_008_),
    .B1(_084_),
    .B2(net27),
    .C1(net34),
    .C2(_010_),
    .ZN(_085_));
 AOI221_X2 _312_ (.A(_080_),
    .B1(_082_),
    .B2(_085_),
    .C1(_041_),
    .C2(_052_),
    .ZN(_086_));
 NAND2_X1 _313_ (.A1(_039_),
    .A2(_081_),
    .ZN(_087_));
 OAI22_X2 _314_ (.A1(_046_),
    .A2(_048_),
    .B1(_087_),
    .B2(_033_),
    .ZN(_088_));
 OAI21_X1 _315_ (.A(_074_),
    .B1(_086_),
    .B2(_088_),
    .ZN(_089_));
 INV_X1 _316_ (.A(net9),
    .ZN(_090_));
 NOR4_X4 _317_ (.A1(_118_),
    .A2(_122_),
    .A3(_119_),
    .A4(_123_),
    .ZN(_091_));
 NOR2_X2 _318_ (.A1(_090_),
    .A2(_091_),
    .ZN(_006_));
 AND3_X1 _319_ (.A1(_064_),
    .A2(_089_),
    .A3(_006_),
    .ZN(_000_));
 NAND3_X2 _320_ (.A1(_135_),
    .A2(_061_),
    .A3(_062_),
    .ZN(_092_));
 NOR2_X1 _321_ (.A1(_057_),
    .A2(_059_),
    .ZN(_093_));
 AOI21_X1 _322_ (.A(_093_),
    .B1(_052_),
    .B2(_041_),
    .ZN(_094_));
 OAI21_X1 _323_ (.A(_010_),
    .B1(_046_),
    .B2(_048_),
    .ZN(_095_));
 OAI221_X2 _324_ (.A(_092_),
    .B1(_051_),
    .B2(_034_),
    .C1(_094_),
    .C2(_095_),
    .ZN(_096_));
 AND3_X1 _325_ (.A1(_096_),
    .A2(_089_),
    .A3(_006_),
    .ZN(_001_));
 OAI211_X2 _326_ (.A(_074_),
    .B(_006_),
    .C1(_088_),
    .C2(_086_),
    .ZN(_097_));
 NOR2_X1 _327_ (.A1(_097_),
    .A2(_096_),
    .ZN(_002_));
 NOR2_X1 _328_ (.A1(_064_),
    .A2(_097_),
    .ZN(_003_));
 NAND2_X1 _329_ (.A1(_126_),
    .A2(_091_),
    .ZN(_098_));
 AOI21_X1 _330_ (.A(_090_),
    .B1(net22),
    .B2(_098_),
    .ZN(_004_));
 NAND2_X1 _331_ (.A1(net15),
    .A2(_091_),
    .ZN(_099_));
 AOI21_X1 _332_ (.A(_090_),
    .B1(_089_),
    .B2(_099_),
    .ZN(_005_));
 HA_X1 _333_ (.A(_142_),
    .B(_143_),
    .CO(_144_),
    .S(_145_));
 HA_X1 _334_ (.A(_146_),
    .B(_147_),
    .CO(_148_),
    .S(_149_));
 HA_X1 _335_ (.A(_150_),
    .B(_151_),
    .CO(_152_),
    .S(_153_));
 HA_X1 _336_ (.A(net33),
    .B(net31),
    .CO(_154_),
    .S(_155_));
 HA_X1 _337_ (.A(net32),
    .B(net15),
    .CO(_156_),
    .S(_157_));
 HA_X1 _338_ (.A(net32),
    .B(net15),
    .CO(_158_),
    .S(_159_));
 HA_X1 _339_ (.A(net14),
    .B(net29),
    .CO(_160_),
    .S(_161_));
 HA_X1 _340_ (.A(net14),
    .B(net30),
    .CO(_162_),
    .S(_163_));
 HA_X1 _341_ (.A(net14),
    .B(net15),
    .CO(_164_),
    .S(_165_));
 HA_X1 _342_ (.A(net14),
    .B(net15),
    .CO(_166_),
    .S(_167_));
 HA_X1 _343_ (.A(_168_),
    .B(_169_),
    .CO(_170_),
    .S(_171_));
 HA_X1 _344_ (.A(_172_),
    .B(_173_),
    .CO(_174_),
    .S(_175_));
 HA_X1 _345_ (.A(_177_),
    .B(_176_),
    .CO(_178_),
    .S(_179_));
 HA_X1 _346_ (.A(_180_),
    .B(_181_),
    .CO(_182_),
    .S(_183_));
 DFF_X1 \grant[0]$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_141_));
 DFF_X1 \grant[1]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_140_));
 DFF_X1 \grant[2]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net12),
    .QN(_139_));
 DFF_X1 \grant[3]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_138_));
 DFF_X2 \last_grant_idx[0]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_150_));
 DFF_X2 \last_grant_idx[1]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net15),
    .QN(_151_));
 DFF_X1 \valid$_SDFF_PN0_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_137_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_57 ();
 BUF_X1 input1 (.A(priorities[0]),
    .Z(net1));
 BUF_X1 input2 (.A(priorities[1]),
    .Z(net2));
 BUF_X2 input3 (.A(priorities[2]),
    .Z(net3));
 BUF_X2 input4 (.A(priorities[3]),
    .Z(net4));
 BUF_X2 input5 (.A(priorities[4]),
    .Z(net5));
 BUF_X2 input6 (.A(priorities[5]),
    .Z(net6));
 BUF_X2 input7 (.A(priorities[6]),
    .Z(net7));
 BUF_X2 input8 (.A(priorities[7]),
    .Z(net8));
 BUF_X1 input9 (.A(rst_n),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(grant[0]));
 BUF_X1 output11 (.A(net11),
    .Z(grant[1]));
 BUF_X1 output12 (.A(net12),
    .Z(grant[2]));
 BUF_X1 output13 (.A(net13),
    .Z(grant[3]));
 BUF_X1 output14 (.A(net14),
    .Z(grant_idx[0]));
 BUF_X1 output15 (.A(net15),
    .Z(grant_idx[1]));
 BUF_X1 output16 (.A(net16),
    .Z(valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 BUF_X2 rebuffer1 (.A(_171_),
    .Z(net17));
 BUF_X1 rebuffer2 (.A(_153_),
    .Z(net18));
 BUF_X1 rebuffer3 (.A(net18),
    .Z(net19));
 BUF_X2 rebuffer4 (.A(_145_),
    .Z(net20));
 BUF_X1 rebuffer5 (.A(net20),
    .Z(net21));
 BUF_X2 rebuffer6 (.A(_064_),
    .Z(net22));
 BUF_X1 rebuffer7 (.A(_124_),
    .Z(net23));
 BUF_X1 rebuffer8 (.A(_124_),
    .Z(net24));
 BUF_X1 rebuffer9 (.A(net24),
    .Z(net25));
 BUF_X1 rebuffer10 (.A(net24),
    .Z(net26));
 BUF_X1 rebuffer11 (.A(_124_),
    .Z(net27));
 BUF_X1 rebuffer12 (.A(net27),
    .Z(net28));
 BUF_X1 rebuffer13 (.A(_151_),
    .Z(net29));
 BUF_X1 rebuffer14 (.A(_151_),
    .Z(net30));
 BUF_X1 rebuffer15 (.A(net30),
    .Z(net31));
 BUF_X1 rebuffer16 (.A(_150_),
    .Z(net32));
 BUF_X1 rebuffer17 (.A(net32),
    .Z(net33));
 BUF_X1 rebuffer18 (.A(_125_),
    .Z(net34));
 BUF_X2 rebuffer19 (.A(net34),
    .Z(net35));
 BUF_X1 rebuffer20 (.A(net35),
    .Z(net36));
 BUF_X1 rebuffer21 (.A(_120_),
    .Z(net37));
 BUF_X1 rebuffer22 (.A(_120_),
    .Z(net38));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X2 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_67 ();
 FILLCELL_X4 FILLER_0_82 ();
 FILLCELL_X2 FILLER_0_102 ();
 FILLCELL_X4 FILLER_0_112 ();
 FILLCELL_X1 FILLER_0_116 ();
 FILLCELL_X2 FILLER_0_120 ();
 FILLCELL_X1 FILLER_0_122 ();
 FILLCELL_X32 FILLER_0_126 ();
 FILLCELL_X32 FILLER_0_158 ();
 FILLCELL_X16 FILLER_0_190 ();
 FILLCELL_X8 FILLER_0_206 ();
 FILLCELL_X4 FILLER_0_214 ();
 FILLCELL_X2 FILLER_0_218 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_41 ();
 FILLCELL_X2 FILLER_1_45 ();
 FILLCELL_X1 FILLER_1_67 ();
 FILLCELL_X32 FILLER_1_110 ();
 FILLCELL_X32 FILLER_1_142 ();
 FILLCELL_X32 FILLER_1_174 ();
 FILLCELL_X8 FILLER_1_206 ();
 FILLCELL_X4 FILLER_1_214 ();
 FILLCELL_X2 FILLER_1_218 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_49 ();
 FILLCELL_X4 FILLER_2_61 ();
 FILLCELL_X4 FILLER_2_79 ();
 FILLCELL_X2 FILLER_2_83 ();
 FILLCELL_X8 FILLER_2_115 ();
 FILLCELL_X1 FILLER_2_123 ();
 FILLCELL_X32 FILLER_2_126 ();
 FILLCELL_X32 FILLER_2_158 ();
 FILLCELL_X16 FILLER_2_190 ();
 FILLCELL_X8 FILLER_2_206 ();
 FILLCELL_X4 FILLER_2_214 ();
 FILLCELL_X2 FILLER_2_218 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X16 FILLER_3_35 ();
 FILLCELL_X4 FILLER_3_51 ();
 FILLCELL_X16 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_81 ();
 FILLCELL_X2 FILLER_3_89 ();
 FILLCELL_X1 FILLER_3_91 ();
 FILLCELL_X2 FILLER_3_106 ();
 FILLCELL_X4 FILLER_3_110 ();
 FILLCELL_X32 FILLER_3_128 ();
 FILLCELL_X32 FILLER_3_160 ();
 FILLCELL_X16 FILLER_3_192 ();
 FILLCELL_X8 FILLER_3_208 ();
 FILLCELL_X4 FILLER_3_216 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X2 FILLER_4_49 ();
 FILLCELL_X1 FILLER_4_64 ();
 FILLCELL_X8 FILLER_4_70 ();
 FILLCELL_X2 FILLER_4_78 ();
 FILLCELL_X8 FILLER_4_82 ();
 FILLCELL_X1 FILLER_4_90 ();
 FILLCELL_X32 FILLER_4_95 ();
 FILLCELL_X32 FILLER_4_127 ();
 FILLCELL_X32 FILLER_4_159 ();
 FILLCELL_X16 FILLER_4_191 ();
 FILLCELL_X8 FILLER_4_207 ();
 FILLCELL_X4 FILLER_4_215 ();
 FILLCELL_X1 FILLER_4_219 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_49 ();
 FILLCELL_X4 FILLER_5_66 ();
 FILLCELL_X2 FILLER_5_70 ();
 FILLCELL_X1 FILLER_5_72 ();
 FILLCELL_X4 FILLER_5_87 ();
 FILLCELL_X8 FILLER_5_98 ();
 FILLCELL_X2 FILLER_5_106 ();
 FILLCELL_X32 FILLER_5_115 ();
 FILLCELL_X32 FILLER_5_147 ();
 FILLCELL_X32 FILLER_5_179 ();
 FILLCELL_X8 FILLER_5_211 ();
 FILLCELL_X1 FILLER_5_219 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_73 ();
 FILLCELL_X2 FILLER_6_77 ();
 FILLCELL_X1 FILLER_6_79 ();
 FILLCELL_X32 FILLER_6_83 ();
 FILLCELL_X4 FILLER_6_115 ();
 FILLCELL_X2 FILLER_6_119 ();
 FILLCELL_X4 FILLER_6_125 ();
 FILLCELL_X1 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_140 ();
 FILLCELL_X32 FILLER_6_172 ();
 FILLCELL_X16 FILLER_6_204 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_17 ();
 FILLCELL_X2 FILLER_7_21 ();
 FILLCELL_X1 FILLER_7_23 ();
 FILLCELL_X8 FILLER_7_44 ();
 FILLCELL_X2 FILLER_7_52 ();
 FILLCELL_X1 FILLER_7_54 ();
 FILLCELL_X2 FILLER_7_68 ();
 FILLCELL_X1 FILLER_7_70 ();
 FILLCELL_X2 FILLER_7_76 ();
 FILLCELL_X2 FILLER_7_89 ();
 FILLCELL_X8 FILLER_7_100 ();
 FILLCELL_X4 FILLER_7_108 ();
 FILLCELL_X2 FILLER_7_112 ();
 FILLCELL_X32 FILLER_7_140 ();
 FILLCELL_X32 FILLER_7_172 ();
 FILLCELL_X16 FILLER_7_204 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_49 ();
 FILLCELL_X2 FILLER_8_53 ();
 FILLCELL_X8 FILLER_8_58 ();
 FILLCELL_X4 FILLER_8_66 ();
 FILLCELL_X2 FILLER_8_70 ();
 FILLCELL_X16 FILLER_8_101 ();
 FILLCELL_X4 FILLER_8_124 ();
 FILLCELL_X2 FILLER_8_128 ();
 FILLCELL_X32 FILLER_8_147 ();
 FILLCELL_X32 FILLER_8_179 ();
 FILLCELL_X8 FILLER_8_211 ();
 FILLCELL_X1 FILLER_8_219 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X2 FILLER_9_85 ();
 FILLCELL_X1 FILLER_9_87 ();
 FILLCELL_X1 FILLER_9_98 ();
 FILLCELL_X16 FILLER_9_103 ();
 FILLCELL_X2 FILLER_9_119 ();
 FILLCELL_X32 FILLER_9_131 ();
 FILLCELL_X32 FILLER_9_163 ();
 FILLCELL_X16 FILLER_9_195 ();
 FILLCELL_X8 FILLER_9_211 ();
 FILLCELL_X1 FILLER_9_219 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_9 ();
 FILLCELL_X32 FILLER_10_51 ();
 FILLCELL_X2 FILLER_10_83 ();
 FILLCELL_X1 FILLER_10_85 ();
 FILLCELL_X1 FILLER_10_97 ();
 FILLCELL_X8 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_121 ();
 FILLCELL_X32 FILLER_10_132 ();
 FILLCELL_X32 FILLER_10_164 ();
 FILLCELL_X16 FILLER_10_196 ();
 FILLCELL_X8 FILLER_10_212 ();
 FILLCELL_X1 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_5 ();
 FILLCELL_X2 FILLER_11_37 ();
 FILLCELL_X1 FILLER_11_39 ();
 FILLCELL_X16 FILLER_11_47 ();
 FILLCELL_X8 FILLER_11_63 ();
 FILLCELL_X8 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_86 ();
 FILLCELL_X1 FILLER_11_88 ();
 FILLCELL_X16 FILLER_11_98 ();
 FILLCELL_X8 FILLER_11_114 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X16 FILLER_11_193 ();
 FILLCELL_X8 FILLER_11_209 ();
 FILLCELL_X2 FILLER_11_217 ();
 FILLCELL_X1 FILLER_11_219 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_33 ();
 FILLCELL_X1 FILLER_12_37 ();
 FILLCELL_X4 FILLER_12_55 ();
 FILLCELL_X2 FILLER_12_59 ();
 FILLCELL_X4 FILLER_12_70 ();
 FILLCELL_X2 FILLER_12_74 ();
 FILLCELL_X1 FILLER_12_79 ();
 FILLCELL_X8 FILLER_12_86 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X32 FILLER_12_128 ();
 FILLCELL_X32 FILLER_12_160 ();
 FILLCELL_X16 FILLER_12_192 ();
 FILLCELL_X8 FILLER_12_208 ();
 FILLCELL_X4 FILLER_12_216 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_20 ();
 FILLCELL_X2 FILLER_13_24 ();
 FILLCELL_X1 FILLER_13_26 ();
 FILLCELL_X2 FILLER_13_30 ();
 FILLCELL_X1 FILLER_13_32 ();
 FILLCELL_X4 FILLER_13_44 ();
 FILLCELL_X1 FILLER_13_48 ();
 FILLCELL_X32 FILLER_13_113 ();
 FILLCELL_X32 FILLER_13_145 ();
 FILLCELL_X32 FILLER_13_177 ();
 FILLCELL_X8 FILLER_13_209 ();
 FILLCELL_X2 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_219 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_16 ();
 FILLCELL_X4 FILLER_14_20 ();
 FILLCELL_X1 FILLER_14_24 ();
 FILLCELL_X16 FILLER_14_38 ();
 FILLCELL_X2 FILLER_14_54 ();
 FILLCELL_X1 FILLER_14_56 ();
 FILLCELL_X2 FILLER_14_67 ();
 FILLCELL_X2 FILLER_14_72 ();
 FILLCELL_X1 FILLER_14_100 ();
 FILLCELL_X1 FILLER_14_104 ();
 FILLCELL_X32 FILLER_14_113 ();
 FILLCELL_X32 FILLER_14_145 ();
 FILLCELL_X32 FILLER_14_177 ();
 FILLCELL_X8 FILLER_14_209 ();
 FILLCELL_X2 FILLER_14_217 ();
 FILLCELL_X1 FILLER_14_219 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X4 FILLER_15_25 ();
 FILLCELL_X1 FILLER_15_29 ();
 FILLCELL_X16 FILLER_15_39 ();
 FILLCELL_X2 FILLER_15_55 ();
 FILLCELL_X2 FILLER_15_79 ();
 FILLCELL_X1 FILLER_15_84 ();
 FILLCELL_X4 FILLER_15_96 ();
 FILLCELL_X4 FILLER_15_102 ();
 FILLCELL_X2 FILLER_15_106 ();
 FILLCELL_X32 FILLER_15_125 ();
 FILLCELL_X32 FILLER_15_157 ();
 FILLCELL_X16 FILLER_15_189 ();
 FILLCELL_X8 FILLER_15_205 ();
 FILLCELL_X4 FILLER_15_213 ();
 FILLCELL_X2 FILLER_15_217 ();
 FILLCELL_X1 FILLER_15_219 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_13 ();
 FILLCELL_X8 FILLER_16_18 ();
 FILLCELL_X2 FILLER_16_26 ();
 FILLCELL_X16 FILLER_16_45 ();
 FILLCELL_X4 FILLER_16_84 ();
 FILLCELL_X2 FILLER_16_88 ();
 FILLCELL_X1 FILLER_16_90 ();
 FILLCELL_X8 FILLER_16_101 ();
 FILLCELL_X2 FILLER_16_109 ();
 FILLCELL_X32 FILLER_16_128 ();
 FILLCELL_X32 FILLER_16_160 ();
 FILLCELL_X16 FILLER_16_192 ();
 FILLCELL_X8 FILLER_16_208 ();
 FILLCELL_X4 FILLER_16_216 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X4 FILLER_17_25 ();
 FILLCELL_X2 FILLER_17_29 ();
 FILLCELL_X32 FILLER_17_36 ();
 FILLCELL_X16 FILLER_17_68 ();
 FILLCELL_X4 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_121 ();
 FILLCELL_X32 FILLER_17_153 ();
 FILLCELL_X32 FILLER_17_185 ();
 FILLCELL_X2 FILLER_17_217 ();
 FILLCELL_X1 FILLER_17_219 ();
 FILLCELL_X8 FILLER_18_9 ();
 FILLCELL_X16 FILLER_18_39 ();
 FILLCELL_X8 FILLER_18_55 ();
 FILLCELL_X1 FILLER_18_63 ();
 FILLCELL_X8 FILLER_18_68 ();
 FILLCELL_X4 FILLER_18_76 ();
 FILLCELL_X8 FILLER_18_98 ();
 FILLCELL_X2 FILLER_18_106 ();
 FILLCELL_X32 FILLER_18_127 ();
 FILLCELL_X32 FILLER_18_159 ();
 FILLCELL_X16 FILLER_18_191 ();
 FILLCELL_X8 FILLER_18_207 ();
 FILLCELL_X4 FILLER_18_215 ();
 FILLCELL_X1 FILLER_18_219 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X8 FILLER_19_10 ();
 FILLCELL_X1 FILLER_19_18 ();
 FILLCELL_X8 FILLER_19_49 ();
 FILLCELL_X2 FILLER_19_57 ();
 FILLCELL_X1 FILLER_19_59 ();
 FILLCELL_X4 FILLER_19_71 ();
 FILLCELL_X2 FILLER_19_75 ();
 FILLCELL_X8 FILLER_19_90 ();
 FILLCELL_X2 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_100 ();
 FILLCELL_X1 FILLER_19_110 ();
 FILLCELL_X32 FILLER_19_120 ();
 FILLCELL_X32 FILLER_19_152 ();
 FILLCELL_X32 FILLER_19_184 ();
 FILLCELL_X4 FILLER_19_216 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X16 FILLER_20_39 ();
 FILLCELL_X4 FILLER_20_55 ();
 FILLCELL_X2 FILLER_20_59 ();
 FILLCELL_X1 FILLER_20_61 ();
 FILLCELL_X16 FILLER_20_66 ();
 FILLCELL_X4 FILLER_20_82 ();
 FILLCELL_X2 FILLER_20_86 ();
 FILLCELL_X1 FILLER_20_88 ();
 FILLCELL_X8 FILLER_20_91 ();
 FILLCELL_X4 FILLER_20_99 ();
 FILLCELL_X2 FILLER_20_103 ();
 FILLCELL_X32 FILLER_20_123 ();
 FILLCELL_X32 FILLER_20_155 ();
 FILLCELL_X32 FILLER_20_187 ();
 FILLCELL_X1 FILLER_20_219 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_9 ();
 FILLCELL_X1 FILLER_21_11 ();
 FILLCELL_X4 FILLER_21_32 ();
 FILLCELL_X2 FILLER_21_36 ();
 FILLCELL_X1 FILLER_21_38 ();
 FILLCELL_X4 FILLER_21_56 ();
 FILLCELL_X4 FILLER_21_64 ();
 FILLCELL_X1 FILLER_21_68 ();
 FILLCELL_X1 FILLER_21_74 ();
 FILLCELL_X8 FILLER_21_77 ();
 FILLCELL_X2 FILLER_21_85 ();
 FILLCELL_X8 FILLER_21_103 ();
 FILLCELL_X2 FILLER_21_111 ();
 FILLCELL_X1 FILLER_21_113 ();
 FILLCELL_X32 FILLER_21_125 ();
 FILLCELL_X32 FILLER_21_157 ();
 FILLCELL_X16 FILLER_21_189 ();
 FILLCELL_X8 FILLER_21_205 ();
 FILLCELL_X4 FILLER_21_213 ();
 FILLCELL_X2 FILLER_21_217 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_17 ();
 FILLCELL_X4 FILLER_22_25 ();
 FILLCELL_X16 FILLER_22_34 ();
 FILLCELL_X8 FILLER_22_50 ();
 FILLCELL_X1 FILLER_22_58 ();
 FILLCELL_X1 FILLER_22_68 ();
 FILLCELL_X2 FILLER_22_75 ();
 FILLCELL_X8 FILLER_22_95 ();
 FILLCELL_X4 FILLER_22_103 ();
 FILLCELL_X2 FILLER_22_115 ();
 FILLCELL_X32 FILLER_22_137 ();
 FILLCELL_X32 FILLER_22_169 ();
 FILLCELL_X16 FILLER_22_201 ();
 FILLCELL_X2 FILLER_22_217 ();
 FILLCELL_X1 FILLER_22_219 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X16 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_49 ();
 FILLCELL_X2 FILLER_23_57 ();
 FILLCELL_X1 FILLER_23_59 ();
 FILLCELL_X1 FILLER_23_64 ();
 FILLCELL_X2 FILLER_23_69 ();
 FILLCELL_X1 FILLER_23_71 ();
 FILLCELL_X32 FILLER_23_93 ();
 FILLCELL_X32 FILLER_23_125 ();
 FILLCELL_X32 FILLER_23_157 ();
 FILLCELL_X16 FILLER_23_189 ();
 FILLCELL_X8 FILLER_23_205 ();
 FILLCELL_X4 FILLER_23_213 ();
 FILLCELL_X2 FILLER_23_217 ();
 FILLCELL_X1 FILLER_23_219 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_50 ();
 FILLCELL_X32 FILLER_24_82 ();
 FILLCELL_X32 FILLER_24_114 ();
 FILLCELL_X32 FILLER_24_146 ();
 FILLCELL_X32 FILLER_24_178 ();
 FILLCELL_X8 FILLER_24_210 ();
 FILLCELL_X2 FILLER_24_218 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X8 FILLER_25_209 ();
 FILLCELL_X2 FILLER_25_217 ();
 FILLCELL_X1 FILLER_25_219 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X16 FILLER_26_65 ();
 FILLCELL_X1 FILLER_26_81 ();
 FILLCELL_X32 FILLER_26_87 ();
 FILLCELL_X32 FILLER_26_119 ();
 FILLCELL_X32 FILLER_26_151 ();
 FILLCELL_X32 FILLER_26_183 ();
 FILLCELL_X4 FILLER_26_215 ();
 FILLCELL_X1 FILLER_26_219 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X16 FILLER_27_193 ();
 FILLCELL_X8 FILLER_27_209 ();
 FILLCELL_X2 FILLER_27_217 ();
 FILLCELL_X1 FILLER_27_219 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X16 FILLER_28_33 ();
 FILLCELL_X16 FILLER_28_52 ();
 FILLCELL_X8 FILLER_28_68 ();
 FILLCELL_X4 FILLER_28_76 ();
 FILLCELL_X2 FILLER_28_80 ();
 FILLCELL_X8 FILLER_28_89 ();
 FILLCELL_X32 FILLER_28_104 ();
 FILLCELL_X32 FILLER_28_136 ();
 FILLCELL_X32 FILLER_28_168 ();
 FILLCELL_X16 FILLER_28_200 ();
 FILLCELL_X4 FILLER_28_216 ();
endmodule
