module jtag_controller (clk,
    dr_shift_en,
    rst_n,
    tck,
    tdi,
    tdo,
    tms,
    trst_n,
    update_dr,
    dr_in,
    dr_out,
    instruction);
 input clk;
 output dr_shift_en;
 input rst_n;
 input tck;
 input tdi;
 output tdo;
 input tms;
 input trst_n;
 output update_dr;
 input [31:0] dr_in;
 output [31:0] dr_out;
 output [4:0] instruction;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire \dr_shift_reg[0] ;
 wire \dr_shift_reg[10] ;
 wire \dr_shift_reg[11] ;
 wire \dr_shift_reg[12] ;
 wire \dr_shift_reg[13] ;
 wire \dr_shift_reg[14] ;
 wire \dr_shift_reg[15] ;
 wire \dr_shift_reg[16] ;
 wire \dr_shift_reg[17] ;
 wire \dr_shift_reg[18] ;
 wire \dr_shift_reg[19] ;
 wire \dr_shift_reg[1] ;
 wire \dr_shift_reg[20] ;
 wire \dr_shift_reg[21] ;
 wire \dr_shift_reg[22] ;
 wire \dr_shift_reg[23] ;
 wire \dr_shift_reg[24] ;
 wire \dr_shift_reg[25] ;
 wire \dr_shift_reg[26] ;
 wire \dr_shift_reg[27] ;
 wire \dr_shift_reg[28] ;
 wire \dr_shift_reg[29] ;
 wire \dr_shift_reg[2] ;
 wire \dr_shift_reg[30] ;
 wire \dr_shift_reg[31] ;
 wire \dr_shift_reg[3] ;
 wire \dr_shift_reg[4] ;
 wire \dr_shift_reg[5] ;
 wire \dr_shift_reg[6] ;
 wire \dr_shift_reg[7] ;
 wire \dr_shift_reg[8] ;
 wire \dr_shift_reg[9] ;
 wire \ir_shift_reg[0] ;
 wire \ir_shift_reg[1] ;
 wire \ir_shift_reg[2] ;
 wire \ir_shift_reg[3] ;
 wire \ir_shift_reg[4] ;
 wire \next_tap_state[0] ;
 wire \next_tap_state[1] ;
 wire \next_tap_state[2] ;
 wire \next_tap_state[3] ;
 wire \tap_state[0] ;
 wire \tap_state[1] ;
 wire \tap_state[2] ;
 wire \tap_state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;

 sky130_fd_sc_hd__clkbuf_4 _202_ (.A(\tap_state[0] ),
    .X(_076_));
 sky130_fd_sc_hd__buf_4 _203_ (.A(\tap_state[2] ),
    .X(_077_));
 sky130_fd_sc_hd__inv_1 _204_ (.A(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor4_4 _205_ (.A(\tap_state[1] ),
    .B(_076_),
    .C(\tap_state[3] ),
    .D(_078_),
    .Y(net69));
 sky130_fd_sc_hd__nand2_1 _206_ (.A(\tap_state[1] ),
    .B(_076_),
    .Y(_079_));
 sky130_fd_sc_hd__buf_2 _207_ (.A(\tap_state[3] ),
    .X(_080_));
 sky130_fd_sc_hd__nor2b_1 _208_ (.A(_077_),
    .B_N(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__nand2_1 _209_ (.A(\ir_shift_reg[0] ),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(\dr_shift_reg[0] ),
    .B(net69),
    .Y(_083_));
 sky130_fd_sc_hd__o21ai_0 _211_ (.A1(_079_),
    .A2(_082_),
    .B1(_083_),
    .Y(_000_));
 sky130_fd_sc_hd__clkinv_2 _212_ (.A(\tap_state[3] ),
    .Y(_084_));
 sky130_fd_sc_hd__nor4_4 _213_ (.A(\tap_state[1] ),
    .B(_076_),
    .C(_084_),
    .D(_077_),
    .Y(_085_));
 sky130_fd_sc_hd__buf_6 _214_ (.A(_085_),
    .X(net76));
 sky130_fd_sc_hd__inv_1 _215_ (.A(net33),
    .Y(_001_));
 sky130_fd_sc_hd__mux2_1 _216_ (.A0(net52),
    .A1(\dr_shift_reg[23] ),
    .S(net76),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _217_ (.A0(net53),
    .A1(\dr_shift_reg[24] ),
    .S(net76),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _218_ (.A0(net54),
    .A1(\dr_shift_reg[25] ),
    .S(net76),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _219_ (.A0(net55),
    .A1(\dr_shift_reg[26] ),
    .S(net76),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _220_ (.A0(net56),
    .A1(\dr_shift_reg[27] ),
    .S(net76),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(net57),
    .A1(\dr_shift_reg[28] ),
    .S(net76),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _222_ (.A0(net58),
    .A1(\dr_shift_reg[29] ),
    .S(net76),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _223_ (.A0(net59),
    .A1(\dr_shift_reg[2] ),
    .S(net76),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _224_ (.A0(net60),
    .A1(\dr_shift_reg[30] ),
    .S(net76),
    .X(_010_));
 sky130_fd_sc_hd__buf_6 _225_ (.A(_085_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _226_ (.A0(net61),
    .A1(\dr_shift_reg[31] ),
    .S(_086_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _227_ (.A0(net62),
    .A1(\dr_shift_reg[3] ),
    .S(_086_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _228_ (.A0(net63),
    .A1(\dr_shift_reg[4] ),
    .S(_086_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _229_ (.A0(net64),
    .A1(\dr_shift_reg[5] ),
    .S(_086_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(net65),
    .A1(\dr_shift_reg[6] ),
    .S(_086_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _231_ (.A0(net66),
    .A1(\dr_shift_reg[7] ),
    .S(_086_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _232_ (.A0(net67),
    .A1(\dr_shift_reg[8] ),
    .S(_086_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _233_ (.A0(net68),
    .A1(\dr_shift_reg[9] ),
    .S(_086_),
    .X(_018_));
 sky130_fd_sc_hd__nor3_4 _234_ (.A(\tap_state[3] ),
    .B(_077_),
    .C(_079_),
    .Y(_087_));
 sky130_fd_sc_hd__buf_6 _235_ (.A(_087_),
    .X(_088_));
 sky130_fd_sc_hd__mux2i_1 _236_ (.A0(\dr_shift_reg[0] ),
    .A1(\dr_shift_reg[1] ),
    .S(net69),
    .Y(_089_));
 sky130_fd_sc_hd__nand2_1 _237_ (.A(net1),
    .B(_088_),
    .Y(_090_));
 sky130_fd_sc_hd__o21ai_0 _238_ (.A1(_088_),
    .A2(_089_),
    .B1(_090_),
    .Y(_019_));
 sky130_fd_sc_hd__or3b_1 _239_ (.A(\tap_state[1] ),
    .B(_076_),
    .C_N(_077_),
    .X(_091_));
 sky130_fd_sc_hd__nand3b_1 _240_ (.A_N(_077_),
    .B(_076_),
    .C(\tap_state[1] ),
    .Y(_092_));
 sky130_fd_sc_hd__a21oi_2 _241_ (.A1(_091_),
    .A2(_092_),
    .B1(_080_),
    .Y(_093_));
 sky130_fd_sc_hd__clkbuf_4 _242_ (.A(_093_),
    .X(_094_));
 sky130_fd_sc_hd__mux2i_1 _243_ (.A0(\dr_shift_reg[11] ),
    .A1(net2),
    .S(_088_),
    .Y(_095_));
 sky130_fd_sc_hd__clkbuf_4 _244_ (.A(_093_),
    .X(_096_));
 sky130_fd_sc_hd__nor2_1 _245_ (.A(\dr_shift_reg[10] ),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__a21oi_1 _246_ (.A1(_094_),
    .A2(_095_),
    .B1(_097_),
    .Y(_020_));
 sky130_fd_sc_hd__mux2i_1 _247_ (.A0(\dr_shift_reg[12] ),
    .A1(net3),
    .S(_088_),
    .Y(_098_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(\dr_shift_reg[11] ),
    .B(_096_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _249_ (.A1(_094_),
    .A2(_098_),
    .B1(_099_),
    .Y(_021_));
 sky130_fd_sc_hd__mux2i_1 _250_ (.A0(\dr_shift_reg[13] ),
    .A1(net4),
    .S(_088_),
    .Y(_100_));
 sky130_fd_sc_hd__nor2_1 _251_ (.A(\dr_shift_reg[12] ),
    .B(_096_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_1 _252_ (.A1(_094_),
    .A2(_100_),
    .B1(_101_),
    .Y(_022_));
 sky130_fd_sc_hd__mux2i_1 _253_ (.A0(\dr_shift_reg[14] ),
    .A1(net5),
    .S(_088_),
    .Y(_102_));
 sky130_fd_sc_hd__nor2_1 _254_ (.A(\dr_shift_reg[13] ),
    .B(_096_),
    .Y(_103_));
 sky130_fd_sc_hd__a21oi_1 _255_ (.A1(_094_),
    .A2(_102_),
    .B1(_103_),
    .Y(_023_));
 sky130_fd_sc_hd__mux2i_1 _256_ (.A0(\dr_shift_reg[15] ),
    .A1(net6),
    .S(_088_),
    .Y(_104_));
 sky130_fd_sc_hd__nor2_1 _257_ (.A(\dr_shift_reg[14] ),
    .B(_096_),
    .Y(_105_));
 sky130_fd_sc_hd__a21oi_1 _258_ (.A1(_094_),
    .A2(_104_),
    .B1(_105_),
    .Y(_024_));
 sky130_fd_sc_hd__mux2i_1 _259_ (.A0(\dr_shift_reg[16] ),
    .A1(net7),
    .S(_088_),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _260_ (.A(\dr_shift_reg[15] ),
    .B(_096_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _261_ (.A1(_094_),
    .A2(_106_),
    .B1(_107_),
    .Y(_025_));
 sky130_fd_sc_hd__buf_6 _262_ (.A(_087_),
    .X(_108_));
 sky130_fd_sc_hd__mux2i_1 _263_ (.A0(\dr_shift_reg[17] ),
    .A1(net8),
    .S(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(\dr_shift_reg[16] ),
    .B(_096_),
    .Y(_110_));
 sky130_fd_sc_hd__a21oi_1 _265_ (.A1(_094_),
    .A2(_109_),
    .B1(_110_),
    .Y(_026_));
 sky130_fd_sc_hd__mux2i_1 _266_ (.A0(\dr_shift_reg[18] ),
    .A1(net9),
    .S(_108_),
    .Y(_111_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(\dr_shift_reg[17] ),
    .B(_096_),
    .Y(_112_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_094_),
    .A2(_111_),
    .B1(_112_),
    .Y(_027_));
 sky130_fd_sc_hd__mux2i_1 _269_ (.A0(\dr_shift_reg[19] ),
    .A1(net10),
    .S(_108_),
    .Y(_113_));
 sky130_fd_sc_hd__nor2_1 _270_ (.A(\dr_shift_reg[18] ),
    .B(_096_),
    .Y(_114_));
 sky130_fd_sc_hd__a21oi_1 _271_ (.A1(_094_),
    .A2(_113_),
    .B1(_114_),
    .Y(_028_));
 sky130_fd_sc_hd__mux2i_1 _272_ (.A0(\dr_shift_reg[20] ),
    .A1(net11),
    .S(_108_),
    .Y(_115_));
 sky130_fd_sc_hd__nor2_1 _273_ (.A(\dr_shift_reg[19] ),
    .B(_096_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_094_),
    .A2(_115_),
    .B1(_116_),
    .Y(_029_));
 sky130_fd_sc_hd__buf_2 _275_ (.A(_093_),
    .X(_117_));
 sky130_fd_sc_hd__mux2i_1 _276_ (.A0(\dr_shift_reg[2] ),
    .A1(net12),
    .S(_108_),
    .Y(_118_));
 sky130_fd_sc_hd__buf_2 _277_ (.A(_093_),
    .X(_119_));
 sky130_fd_sc_hd__nor2_1 _278_ (.A(\dr_shift_reg[1] ),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(_117_),
    .A2(_118_),
    .B1(_120_),
    .Y(_030_));
 sky130_fd_sc_hd__mux2i_1 _280_ (.A0(\dr_shift_reg[21] ),
    .A1(net13),
    .S(_108_),
    .Y(_121_));
 sky130_fd_sc_hd__nor2_1 _281_ (.A(\dr_shift_reg[20] ),
    .B(_119_),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _282_ (.A1(_117_),
    .A2(_121_),
    .B1(_122_),
    .Y(_031_));
 sky130_fd_sc_hd__mux2i_1 _283_ (.A0(\dr_shift_reg[22] ),
    .A1(net14),
    .S(_108_),
    .Y(_123_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(\dr_shift_reg[21] ),
    .B(_119_),
    .Y(_124_));
 sky130_fd_sc_hd__a21oi_1 _285_ (.A1(_117_),
    .A2(_123_),
    .B1(_124_),
    .Y(_032_));
 sky130_fd_sc_hd__mux2i_1 _286_ (.A0(\dr_shift_reg[23] ),
    .A1(net15),
    .S(_108_),
    .Y(_125_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(\dr_shift_reg[22] ),
    .B(_119_),
    .Y(_126_));
 sky130_fd_sc_hd__a21oi_1 _288_ (.A1(_117_),
    .A2(_125_),
    .B1(_126_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2i_1 _289_ (.A0(\dr_shift_reg[24] ),
    .A1(net16),
    .S(_108_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _290_ (.A(\dr_shift_reg[23] ),
    .B(_119_),
    .Y(_128_));
 sky130_fd_sc_hd__a21oi_1 _291_ (.A1(_117_),
    .A2(_127_),
    .B1(_128_),
    .Y(_034_));
 sky130_fd_sc_hd__mux2i_1 _292_ (.A0(\dr_shift_reg[25] ),
    .A1(net17),
    .S(_108_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _293_ (.A(\dr_shift_reg[24] ),
    .B(_119_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_1 _294_ (.A1(_117_),
    .A2(_129_),
    .B1(_130_),
    .Y(_035_));
 sky130_fd_sc_hd__buf_6 _295_ (.A(_087_),
    .X(_131_));
 sky130_fd_sc_hd__mux2i_1 _296_ (.A0(\dr_shift_reg[26] ),
    .A1(net18),
    .S(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2_1 _297_ (.A(\dr_shift_reg[25] ),
    .B(_119_),
    .Y(_133_));
 sky130_fd_sc_hd__a21oi_1 _298_ (.A1(_117_),
    .A2(_132_),
    .B1(_133_),
    .Y(_036_));
 sky130_fd_sc_hd__mux2i_1 _299_ (.A0(\dr_shift_reg[27] ),
    .A1(net19),
    .S(_131_),
    .Y(_134_));
 sky130_fd_sc_hd__nor2_1 _300_ (.A(\dr_shift_reg[26] ),
    .B(_119_),
    .Y(_135_));
 sky130_fd_sc_hd__a21oi_1 _301_ (.A1(_117_),
    .A2(_134_),
    .B1(_135_),
    .Y(_037_));
 sky130_fd_sc_hd__mux2i_1 _302_ (.A0(\dr_shift_reg[28] ),
    .A1(net20),
    .S(_131_),
    .Y(_136_));
 sky130_fd_sc_hd__nor2_1 _303_ (.A(\dr_shift_reg[27] ),
    .B(_119_),
    .Y(_137_));
 sky130_fd_sc_hd__a21oi_1 _304_ (.A1(_117_),
    .A2(_136_),
    .B1(_137_),
    .Y(_038_));
 sky130_fd_sc_hd__mux2i_1 _305_ (.A0(\dr_shift_reg[29] ),
    .A1(net21),
    .S(_131_),
    .Y(_138_));
 sky130_fd_sc_hd__nor2_1 _306_ (.A(\dr_shift_reg[28] ),
    .B(_119_),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_1 _307_ (.A1(_117_),
    .A2(_138_),
    .B1(_139_),
    .Y(_039_));
 sky130_fd_sc_hd__buf_2 _308_ (.A(_093_),
    .X(_140_));
 sky130_fd_sc_hd__mux2i_1 _309_ (.A0(\dr_shift_reg[30] ),
    .A1(net22),
    .S(_131_),
    .Y(_141_));
 sky130_fd_sc_hd__buf_2 _310_ (.A(_093_),
    .X(_142_));
 sky130_fd_sc_hd__nor2_1 _311_ (.A(\dr_shift_reg[29] ),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a21oi_1 _312_ (.A1(_140_),
    .A2(_141_),
    .B1(_143_),
    .Y(_040_));
 sky130_fd_sc_hd__mux2i_1 _313_ (.A0(\dr_shift_reg[3] ),
    .A1(net23),
    .S(_131_),
    .Y(_144_));
 sky130_fd_sc_hd__nor2_1 _314_ (.A(\dr_shift_reg[2] ),
    .B(_142_),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _315_ (.A1(_140_),
    .A2(_144_),
    .B1(_145_),
    .Y(_041_));
 sky130_fd_sc_hd__mux2i_1 _316_ (.A0(\dr_shift_reg[30] ),
    .A1(\dr_shift_reg[31] ),
    .S(net69),
    .Y(_146_));
 sky130_fd_sc_hd__nand2_1 _317_ (.A(net24),
    .B(_088_),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_0 _318_ (.A1(_088_),
    .A2(_146_),
    .B1(_147_),
    .Y(_042_));
 sky130_fd_sc_hd__mux2i_1 _319_ (.A0(net34),
    .A1(net25),
    .S(_131_),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(\dr_shift_reg[31] ),
    .B(_142_),
    .Y(_149_));
 sky130_fd_sc_hd__a21oi_1 _321_ (.A1(_140_),
    .A2(_148_),
    .B1(_149_),
    .Y(_043_));
 sky130_fd_sc_hd__mux2i_1 _322_ (.A0(\dr_shift_reg[4] ),
    .A1(net26),
    .S(_131_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _323_ (.A(\dr_shift_reg[3] ),
    .B(_142_),
    .Y(_151_));
 sky130_fd_sc_hd__a21oi_1 _324_ (.A1(_140_),
    .A2(_150_),
    .B1(_151_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2i_1 _325_ (.A0(\dr_shift_reg[5] ),
    .A1(net27),
    .S(_131_),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_1 _326_ (.A(\dr_shift_reg[4] ),
    .B(_142_),
    .Y(_153_));
 sky130_fd_sc_hd__a21oi_1 _327_ (.A1(_140_),
    .A2(_152_),
    .B1(_153_),
    .Y(_045_));
 sky130_fd_sc_hd__mux2i_1 _328_ (.A0(\dr_shift_reg[6] ),
    .A1(net28),
    .S(_131_),
    .Y(_154_));
 sky130_fd_sc_hd__nor2_1 _329_ (.A(\dr_shift_reg[5] ),
    .B(_142_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_1 _330_ (.A1(_140_),
    .A2(_154_),
    .B1(_155_),
    .Y(_046_));
 sky130_fd_sc_hd__mux2i_1 _331_ (.A0(\dr_shift_reg[7] ),
    .A1(net29),
    .S(_087_),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_1 _332_ (.A(\dr_shift_reg[6] ),
    .B(_142_),
    .Y(_157_));
 sky130_fd_sc_hd__a21oi_1 _333_ (.A1(_140_),
    .A2(_156_),
    .B1(_157_),
    .Y(_047_));
 sky130_fd_sc_hd__mux2i_1 _334_ (.A0(\dr_shift_reg[8] ),
    .A1(net30),
    .S(_087_),
    .Y(_158_));
 sky130_fd_sc_hd__nor2_1 _335_ (.A(\dr_shift_reg[7] ),
    .B(_142_),
    .Y(_159_));
 sky130_fd_sc_hd__a21oi_1 _336_ (.A1(_140_),
    .A2(_158_),
    .B1(_159_),
    .Y(_048_));
 sky130_fd_sc_hd__mux2i_1 _337_ (.A0(\dr_shift_reg[9] ),
    .A1(net31),
    .S(_087_),
    .Y(_160_));
 sky130_fd_sc_hd__nor2_1 _338_ (.A(\dr_shift_reg[8] ),
    .B(_142_),
    .Y(_161_));
 sky130_fd_sc_hd__a21oi_1 _339_ (.A1(_140_),
    .A2(_160_),
    .B1(_161_),
    .Y(_049_));
 sky130_fd_sc_hd__mux2i_1 _340_ (.A0(\dr_shift_reg[10] ),
    .A1(net32),
    .S(_087_),
    .Y(_162_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(\dr_shift_reg[9] ),
    .B(_142_),
    .Y(_163_));
 sky130_fd_sc_hd__a21oi_1 _342_ (.A1(_140_),
    .A2(_162_),
    .B1(_163_),
    .Y(_050_));
 sky130_fd_sc_hd__buf_2 _343_ (.A(\tap_state[1] ),
    .X(_164_));
 sky130_fd_sc_hd__nand2_2 _344_ (.A(_164_),
    .B(_081_),
    .Y(_165_));
 sky130_fd_sc_hd__buf_2 _345_ (.A(_076_),
    .X(_166_));
 sky130_fd_sc_hd__clkinvlp_4 _346_ (.A(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_1 _347_ (.A(_167_),
    .B(\ir_shift_reg[1] ),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(\ir_shift_reg[0] ),
    .B(_165_),
    .Y(_169_));
 sky130_fd_sc_hd__o21ai_0 _349_ (.A1(_165_),
    .A2(_168_),
    .B1(_169_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2_1 _350_ (.A(_167_),
    .B(\ir_shift_reg[2] ),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _351_ (.A(\ir_shift_reg[1] ),
    .B(_165_),
    .Y(_171_));
 sky130_fd_sc_hd__o21ai_0 _352_ (.A1(_165_),
    .A2(_170_),
    .B1(_171_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_1 _353_ (.A(_167_),
    .B(\ir_shift_reg[3] ),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _354_ (.A(\ir_shift_reg[2] ),
    .B(_165_),
    .Y(_173_));
 sky130_fd_sc_hd__o21ai_0 _355_ (.A1(_165_),
    .A2(_172_),
    .B1(_173_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _356_ (.A(_167_),
    .B(\ir_shift_reg[4] ),
    .Y(_174_));
 sky130_fd_sc_hd__nand2_1 _357_ (.A(\ir_shift_reg[3] ),
    .B(_165_),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _358_ (.A1(_165_),
    .A2(_174_),
    .B1(_175_),
    .Y(_059_));
 sky130_fd_sc_hd__nand2_1 _359_ (.A(_166_),
    .B(net34),
    .Y(_176_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(\ir_shift_reg[4] ),
    .B(_165_),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_0 _361_ (.A1(_165_),
    .A2(_176_),
    .B1(_177_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(net37),
    .A1(\dr_shift_reg[0] ),
    .S(_086_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(net38),
    .A1(\dr_shift_reg[10] ),
    .S(_086_),
    .X(_062_));
 sky130_fd_sc_hd__buf_6 _364_ (.A(_085_),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(net39),
    .A1(\dr_shift_reg[11] ),
    .S(_178_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _366_ (.A0(net40),
    .A1(\dr_shift_reg[12] ),
    .S(_178_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(net41),
    .A1(\dr_shift_reg[13] ),
    .S(_178_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _368_ (.A0(net42),
    .A1(\dr_shift_reg[14] ),
    .S(_178_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(net43),
    .A1(\dr_shift_reg[15] ),
    .S(_178_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(net44),
    .A1(\dr_shift_reg[16] ),
    .S(_178_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(net45),
    .A1(\dr_shift_reg[17] ),
    .S(_178_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(net46),
    .A1(\dr_shift_reg[18] ),
    .S(_178_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(net47),
    .A1(\dr_shift_reg[19] ),
    .S(_178_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(net48),
    .A1(\dr_shift_reg[1] ),
    .S(_178_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(net49),
    .A1(\dr_shift_reg[20] ),
    .S(_085_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(net50),
    .A1(\dr_shift_reg[21] ),
    .S(_085_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(net51),
    .A1(\dr_shift_reg[22] ),
    .S(_085_),
    .X(_075_));
 sky130_fd_sc_hd__buf_2 _378_ (.A(_077_),
    .X(_179_));
 sky130_fd_sc_hd__nand4_4 _379_ (.A(_164_),
    .B(_076_),
    .C(_080_),
    .D(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(\ir_shift_reg[0] ),
    .A1(net70),
    .S(_180_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(\ir_shift_reg[1] ),
    .A1(net71),
    .S(_180_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(\ir_shift_reg[2] ),
    .A1(net72),
    .S(_180_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(\ir_shift_reg[3] ),
    .A1(net73),
    .S(_180_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(\ir_shift_reg[4] ),
    .A1(net74),
    .S(_180_),
    .X(_055_));
 sky130_fd_sc_hd__buf_2 _385_ (.A(net35),
    .X(_181_));
 sky130_fd_sc_hd__inv_1 _386_ (.A(net35),
    .Y(_182_));
 sky130_fd_sc_hd__a21oi_1 _387_ (.A1(_164_),
    .A2(_182_),
    .B1(_179_),
    .Y(_183_));
 sky130_fd_sc_hd__o22ai_1 _388_ (.A1(_078_),
    .A2(_181_),
    .B1(_183_),
    .B2(_167_),
    .Y(_184_));
 sky130_fd_sc_hd__a21oi_1 _389_ (.A1(_166_),
    .A2(_080_),
    .B1(_181_),
    .Y(_185_));
 sky130_fd_sc_hd__o211ai_1 _390_ (.A1(_166_),
    .A2(_078_),
    .B1(_181_),
    .C1(_080_),
    .Y(_186_));
 sky130_fd_sc_hd__o31ai_1 _391_ (.A1(_164_),
    .A2(_179_),
    .A3(_185_),
    .B1(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a21oi_1 _392_ (.A1(_084_),
    .A2(_184_),
    .B1(_187_),
    .Y(\next_tap_state[0] ));
 sky130_fd_sc_hd__xnor2_1 _393_ (.A(_179_),
    .B(_181_),
    .Y(_188_));
 sky130_fd_sc_hd__nor3_1 _394_ (.A(_164_),
    .B(_080_),
    .C(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__a21oi_1 _395_ (.A1(_182_),
    .A2(_081_),
    .B1(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__a21oi_1 _396_ (.A1(_080_),
    .A2(_181_),
    .B1(_164_),
    .Y(_191_));
 sky130_fd_sc_hd__a311oi_1 _397_ (.A1(_164_),
    .A2(_078_),
    .A3(_181_),
    .B1(_191_),
    .C1(_166_),
    .Y(_192_));
 sky130_fd_sc_hd__a31oi_1 _398_ (.A1(_080_),
    .A2(_179_),
    .A3(_181_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__o21ai_0 _399_ (.A1(_167_),
    .A2(_190_),
    .B1(_193_),
    .Y(\next_tap_state[1] ));
 sky130_fd_sc_hd__nand3_1 _400_ (.A(_166_),
    .B(_179_),
    .C(_181_),
    .Y(_194_));
 sky130_fd_sc_hd__o21ai_0 _401_ (.A1(_084_),
    .A2(_181_),
    .B1(_194_),
    .Y(_195_));
 sky130_fd_sc_hd__nand3_1 _402_ (.A(_166_),
    .B(_084_),
    .C(_181_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _403_ (.A1(_179_),
    .A2(_196_),
    .B1(_164_),
    .Y(_197_));
 sky130_fd_sc_hd__nor3_1 _404_ (.A(_166_),
    .B(_080_),
    .C(_179_),
    .Y(_198_));
 sky130_fd_sc_hd__a211oi_1 _405_ (.A1(_164_),
    .A2(_195_),
    .B1(_197_),
    .C1(_198_),
    .Y(\next_tap_state[2] ));
 sky130_fd_sc_hd__a21oi_1 _406_ (.A1(_166_),
    .A2(_182_),
    .B1(_164_),
    .Y(_199_));
 sky130_fd_sc_hd__a21oi_1 _407_ (.A1(_166_),
    .A2(_084_),
    .B1(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__a21oi_1 _408_ (.A1(_167_),
    .A2(_179_),
    .B1(_182_),
    .Y(_201_));
 sky130_fd_sc_hd__o221a_1 _409_ (.A1(_179_),
    .A2(_200_),
    .B1(_201_),
    .B2(_080_),
    .C1(_180_),
    .X(\next_tap_state[3] ));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[0]$_DFFE_NN0P_  (.D(_061_),
    .Q(net37),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[10]$_DFFE_NN0P_  (.D(_062_),
    .Q(net38),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[11]$_DFFE_NN0P_  (.D(_063_),
    .Q(net39),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[12]$_DFFE_NN0P_  (.D(_064_),
    .Q(net40),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[13]$_DFFE_NN0P_  (.D(_065_),
    .Q(net41),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[14]$_DFFE_NN0P_  (.D(_066_),
    .Q(net42),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[15]$_DFFE_NN0P_  (.D(_067_),
    .Q(net43),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[16]$_DFFE_NN0P_  (.D(_068_),
    .Q(net44),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[17]$_DFFE_NN0P_  (.D(_069_),
    .Q(net45),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[18]$_DFFE_NN0P_  (.D(_070_),
    .Q(net46),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[19]$_DFFE_NN0P_  (.D(_071_),
    .Q(net47),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[1]$_DFFE_NN0P_  (.D(_072_),
    .Q(net48),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[20]$_DFFE_NN0P_  (.D(_073_),
    .Q(net49),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[21]$_DFFE_NN0P_  (.D(_074_),
    .Q(net50),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[22]$_DFFE_NN0P_  (.D(_075_),
    .Q(net51),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[23]$_DFFE_NN0P_  (.D(_002_),
    .Q(net52),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[24]$_DFFE_NN0P_  (.D(_003_),
    .Q(net53),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[25]$_DFFE_NN0P_  (.D(_004_),
    .Q(net54),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[26]$_DFFE_NN0P_  (.D(_005_),
    .Q(net55),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[27]$_DFFE_NN0P_  (.D(_006_),
    .Q(net56),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[28]$_DFFE_NN0P_  (.D(_007_),
    .Q(net57),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[29]$_DFFE_NN0P_  (.D(_008_),
    .Q(net58),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[2]$_DFFE_NN0P_  (.D(_009_),
    .Q(net59),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[30]$_DFFE_NN0P_  (.D(_010_),
    .Q(net60),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[31]$_DFFE_NN0P_  (.D(_011_),
    .Q(net61),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[3]$_DFFE_NN0P_  (.D(_012_),
    .Q(net62),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[4]$_DFFE_NN0P_  (.D(_013_),
    .Q(net63),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[5]$_DFFE_NN0P_  (.D(_014_),
    .Q(net64),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[6]$_DFFE_NN0P_  (.D(_015_),
    .Q(net65),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[7]$_DFFE_NN0P_  (.D(_016_),
    .Q(net66),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[8]$_DFFE_NN0P_  (.D(_017_),
    .Q(net67),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \dr_reg[9]$_DFFE_NN0P_  (.D(_018_),
    .Q(net68),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[0]$_DFFE_PN0P_  (.D(_019_),
    .Q(\dr_shift_reg[0] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[10]$_DFFE_PN0P_  (.D(_020_),
    .Q(\dr_shift_reg[10] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[11]$_DFFE_PN0P_  (.D(_021_),
    .Q(\dr_shift_reg[11] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[12]$_DFFE_PN0P_  (.D(_022_),
    .Q(\dr_shift_reg[12] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[13]$_DFFE_PN0P_  (.D(_023_),
    .Q(\dr_shift_reg[13] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[14]$_DFFE_PN0P_  (.D(_024_),
    .Q(\dr_shift_reg[14] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[15]$_DFFE_PN0P_  (.D(_025_),
    .Q(\dr_shift_reg[15] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[16]$_DFFE_PN0P_  (.D(_026_),
    .Q(\dr_shift_reg[16] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[17]$_DFFE_PN0P_  (.D(_027_),
    .Q(\dr_shift_reg[17] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[18]$_DFFE_PN0P_  (.D(_028_),
    .Q(\dr_shift_reg[18] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[19]$_DFFE_PN0P_  (.D(_029_),
    .Q(\dr_shift_reg[19] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[1]$_DFFE_PN0P_  (.D(_030_),
    .Q(\dr_shift_reg[1] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[20]$_DFFE_PN0P_  (.D(_031_),
    .Q(\dr_shift_reg[20] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[21]$_DFFE_PN0P_  (.D(_032_),
    .Q(\dr_shift_reg[21] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[22]$_DFFE_PN0P_  (.D(_033_),
    .Q(\dr_shift_reg[22] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[23]$_DFFE_PN0P_  (.D(_034_),
    .Q(\dr_shift_reg[23] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[24]$_DFFE_PN0P_  (.D(_035_),
    .Q(\dr_shift_reg[24] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[25]$_DFFE_PN0P_  (.D(_036_),
    .Q(\dr_shift_reg[25] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[26]$_DFFE_PN0P_  (.D(_037_),
    .Q(\dr_shift_reg[26] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[27]$_DFFE_PN0P_  (.D(_038_),
    .Q(\dr_shift_reg[27] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[28]$_DFFE_PN0P_  (.D(_039_),
    .Q(\dr_shift_reg[28] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[29]$_DFFE_PN0P_  (.D(_040_),
    .Q(\dr_shift_reg[29] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[2]$_DFFE_PN0P_  (.D(_041_),
    .Q(\dr_shift_reg[2] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[30]$_DFFE_PN0P_  (.D(_042_),
    .Q(\dr_shift_reg[30] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[31]$_DFFE_PN0P_  (.D(_043_),
    .Q(\dr_shift_reg[31] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[3]$_DFFE_PN0P_  (.D(_044_),
    .Q(\dr_shift_reg[3] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[4]$_DFFE_PN0P_  (.D(_045_),
    .Q(\dr_shift_reg[4] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[5]$_DFFE_PN0P_  (.D(_046_),
    .Q(\dr_shift_reg[5] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[6]$_DFFE_PN0P_  (.D(_047_),
    .Q(\dr_shift_reg[6] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[7]$_DFFE_PN0P_  (.D(_048_),
    .Q(\dr_shift_reg[7] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[8]$_DFFE_PN0P_  (.D(_049_),
    .Q(\dr_shift_reg[8] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \dr_shift_reg[9]$_DFFE_PN0P_  (.D(_050_),
    .Q(\dr_shift_reg[9] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfstp_1 \ir_reg[0]$_DFFE_NN1N_  (.D(_051_),
    .Q(net70),
    .SET_B(net36),
    .CLK(_001_));
 sky130_fd_sc_hd__dfrtn_1 \ir_reg[1]$_DFFE_NN0N_  (.D(_052_),
    .Q(net71),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \ir_reg[2]$_DFFE_NN0N_  (.D(_053_),
    .Q(net72),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \ir_reg[3]$_DFFE_NN0N_  (.D(_054_),
    .Q(net73),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfrtn_1 \ir_reg[4]$_DFFE_NN0N_  (.D(_055_),
    .Q(net74),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__dfstp_1 \ir_shift_reg[0]$_DFFE_PN1P_  (.D(_056_),
    .Q(\ir_shift_reg[0] ),
    .SET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \ir_shift_reg[1]$_DFFE_PN0P_  (.D(_057_),
    .Q(\ir_shift_reg[1] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \ir_shift_reg[2]$_DFFE_PN0P_  (.D(_058_),
    .Q(\ir_shift_reg[2] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \ir_shift_reg[3]$_DFFE_PN0P_  (.D(_059_),
    .Q(\ir_shift_reg[3] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \ir_shift_reg[4]$_DFFE_PN0P_  (.D(_060_),
    .Q(\ir_shift_reg[4] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \tap_state[0]$_DFF_PN0_  (.D(\next_tap_state[0] ),
    .Q(\tap_state[0] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_4 \tap_state[1]$_DFF_PN0_  (.D(\next_tap_state[1] ),
    .Q(\tap_state[1] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_1 \tap_state[2]$_DFF_PN0_  (.D(\next_tap_state[2] ),
    .Q(\tap_state[2] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtp_2 \tap_state[3]$_DFF_PN0_  (.D(\next_tap_state[3] ),
    .Q(\tap_state[3] ),
    .RESET_B(net36),
    .CLK(net33));
 sky130_fd_sc_hd__dfrtn_1 \tdo_mux$_DFF_NN0_  (.D(_000_),
    .Q(net75),
    .RESET_B(net36),
    .CLK_N(net33));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_74 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(dr_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dr_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(dr_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(dr_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(dr_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(dr_in[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(dr_in[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(dr_in[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(dr_in[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(dr_in[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(dr_in[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(dr_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(dr_in[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(dr_in[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(dr_in[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(dr_in[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(dr_in[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(dr_in[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(dr_in[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(dr_in[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(dr_in[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(dr_in[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(dr_in[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(dr_in[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(dr_in[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(dr_in[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(dr_in[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(dr_in[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(dr_in[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(dr_in[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(dr_in[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(dr_in[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_16 input33 (.A(tck),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(tdi),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(tms),
    .X(net35));
 sky130_fd_sc_hd__buf_16 input36 (.A(trst_n),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(dr_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(dr_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(dr_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(dr_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(dr_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(dr_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(dr_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(dr_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(dr_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(dr_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(dr_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(dr_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(dr_out[20]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(dr_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(dr_out[22]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(dr_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(dr_out[24]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(dr_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(dr_out[26]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(dr_out[27]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(dr_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(dr_out[29]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(dr_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(dr_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(dr_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(dr_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(dr_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(dr_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(dr_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(dr_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(dr_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(dr_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(dr_shift_en));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(instruction[0]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(instruction[1]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(instruction[2]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(instruction[3]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(instruction[4]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(tdo));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(update_dr));
 sky130_fd_sc_hd__fill_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_167 ();
endmodule
