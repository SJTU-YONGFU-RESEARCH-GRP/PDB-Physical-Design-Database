module dma_controller (clk,
    debug_has_active_channels,
    rst_n,
    channel_busy,
    channel_done,
    channel_dst_addr,
    channel_enable,
    channel_error,
    channel_length,
    channel_mode,
    channel_src_addr,
    channel_start,
    debug_active_channels,
    debug_channel_state,
    debug_transfer_count,
    dst_addr,
    dst_wdata,
    dst_wready,
    dst_write,
    dst_wstrb,
    src_addr,
    src_rdata,
    src_read,
    src_rready,
    src_rvalid);
 input clk;
 output debug_has_active_channels;
 input rst_n;
 output [3:0] channel_busy;
 output [3:0] channel_done;
 input [127:0] channel_dst_addr;
 input [3:0] channel_enable;
 output [3:0] channel_error;
 input [127:0] channel_length;
 input [7:0] channel_mode;
 input [127:0] channel_src_addr;
 input [3:0] channel_start;
 output [3:0] debug_active_channels;
 output [11:0] debug_channel_state;
 output [127:0] debug_transfer_count;
 output [127:0] dst_addr;
 output [127:0] dst_wdata;
 input [3:0] dst_wready;
 output [3:0] dst_write;
 output [15:0] dst_wstrb;
 output [127:0] src_addr;
 input [127:0] src_rdata;
 output [3:0] src_read;
 output [3:0] src_rready;
 input [3:0] src_rvalid;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire clknet_0_clk;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire \active_channel_count[0] ;
 wire \active_channel_count[1] ;
 wire \active_channel_count[2] ;
 wire \active_channel_count[3] ;
 wire \channel_state[0][0] ;
 wire \channel_state[0][1] ;
 wire \channel_state[0][2] ;
 wire \channel_state[1][0] ;
 wire \channel_state[1][1] ;
 wire \channel_state[1][2] ;
 wire \channel_state[2][0] ;
 wire \channel_state[2][1] ;
 wire \channel_state[2][2] ;
 wire \channel_state[3][0] ;
 wire \channel_state[3][1] ;
 wire \channel_state[3][2] ;
 wire \transfer_count[0][0] ;
 wire \transfer_count[0][10] ;
 wire \transfer_count[0][11] ;
 wire \transfer_count[0][12] ;
 wire \transfer_count[0][13] ;
 wire \transfer_count[0][14] ;
 wire \transfer_count[0][15] ;
 wire \transfer_count[0][16] ;
 wire \transfer_count[0][17] ;
 wire \transfer_count[0][18] ;
 wire \transfer_count[0][19] ;
 wire \transfer_count[0][1] ;
 wire \transfer_count[0][20] ;
 wire \transfer_count[0][21] ;
 wire \transfer_count[0][22] ;
 wire \transfer_count[0][23] ;
 wire \transfer_count[0][24] ;
 wire \transfer_count[0][25] ;
 wire \transfer_count[0][26] ;
 wire \transfer_count[0][27] ;
 wire \transfer_count[0][28] ;
 wire \transfer_count[0][29] ;
 wire \transfer_count[0][2] ;
 wire \transfer_count[0][30] ;
 wire \transfer_count[0][31] ;
 wire \transfer_count[0][3] ;
 wire \transfer_count[0][4] ;
 wire \transfer_count[0][5] ;
 wire \transfer_count[0][6] ;
 wire \transfer_count[0][7] ;
 wire \transfer_count[0][8] ;
 wire \transfer_count[0][9] ;
 wire \transfer_count[1][0] ;
 wire \transfer_count[1][10] ;
 wire \transfer_count[1][11] ;
 wire \transfer_count[1][12] ;
 wire \transfer_count[1][13] ;
 wire \transfer_count[1][14] ;
 wire \transfer_count[1][15] ;
 wire \transfer_count[1][16] ;
 wire \transfer_count[1][17] ;
 wire \transfer_count[1][18] ;
 wire \transfer_count[1][19] ;
 wire \transfer_count[1][1] ;
 wire \transfer_count[1][20] ;
 wire \transfer_count[1][21] ;
 wire \transfer_count[1][22] ;
 wire \transfer_count[1][23] ;
 wire \transfer_count[1][24] ;
 wire \transfer_count[1][25] ;
 wire \transfer_count[1][26] ;
 wire \transfer_count[1][27] ;
 wire \transfer_count[1][28] ;
 wire \transfer_count[1][29] ;
 wire \transfer_count[1][2] ;
 wire \transfer_count[1][30] ;
 wire \transfer_count[1][31] ;
 wire \transfer_count[1][3] ;
 wire \transfer_count[1][4] ;
 wire \transfer_count[1][5] ;
 wire \transfer_count[1][6] ;
 wire \transfer_count[1][7] ;
 wire \transfer_count[1][8] ;
 wire \transfer_count[1][9] ;
 wire \transfer_count[2][0] ;
 wire \transfer_count[2][10] ;
 wire \transfer_count[2][11] ;
 wire \transfer_count[2][12] ;
 wire \transfer_count[2][13] ;
 wire \transfer_count[2][14] ;
 wire \transfer_count[2][15] ;
 wire \transfer_count[2][16] ;
 wire \transfer_count[2][17] ;
 wire \transfer_count[2][18] ;
 wire \transfer_count[2][19] ;
 wire \transfer_count[2][1] ;
 wire \transfer_count[2][20] ;
 wire \transfer_count[2][21] ;
 wire \transfer_count[2][22] ;
 wire \transfer_count[2][23] ;
 wire \transfer_count[2][24] ;
 wire \transfer_count[2][25] ;
 wire \transfer_count[2][26] ;
 wire \transfer_count[2][27] ;
 wire \transfer_count[2][28] ;
 wire \transfer_count[2][29] ;
 wire \transfer_count[2][2] ;
 wire \transfer_count[2][30] ;
 wire \transfer_count[2][31] ;
 wire \transfer_count[2][3] ;
 wire \transfer_count[2][4] ;
 wire \transfer_count[2][5] ;
 wire \transfer_count[2][6] ;
 wire \transfer_count[2][7] ;
 wire \transfer_count[2][8] ;
 wire \transfer_count[2][9] ;
 wire \transfer_count[3][0] ;
 wire \transfer_count[3][10] ;
 wire \transfer_count[3][11] ;
 wire \transfer_count[3][12] ;
 wire \transfer_count[3][13] ;
 wire \transfer_count[3][14] ;
 wire \transfer_count[3][15] ;
 wire \transfer_count[3][16] ;
 wire \transfer_count[3][17] ;
 wire \transfer_count[3][18] ;
 wire \transfer_count[3][19] ;
 wire \transfer_count[3][1] ;
 wire \transfer_count[3][20] ;
 wire \transfer_count[3][21] ;
 wire \transfer_count[3][22] ;
 wire \transfer_count[3][23] ;
 wire \transfer_count[3][24] ;
 wire \transfer_count[3][25] ;
 wire \transfer_count[3][26] ;
 wire \transfer_count[3][27] ;
 wire \transfer_count[3][28] ;
 wire \transfer_count[3][29] ;
 wire \transfer_count[3][2] ;
 wire \transfer_count[3][30] ;
 wire \transfer_count[3][31] ;
 wire \transfer_count[3][3] ;
 wire \transfer_count[3][4] ;
 wire \transfer_count[3][5] ;
 wire \transfer_count[3][6] ;
 wire \transfer_count[3][7] ;
 wire \transfer_count[3][8] ;
 wire \transfer_count[3][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__nand2_1 _1443_ (.A(\transfer_count[1][2] ),
    .B(\transfer_count[1][3] ),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_2 _1444_ (.A(\transfer_count[1][4] ),
    .B(\transfer_count[1][5] ),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(\transfer_count[1][0] ),
    .B(\transfer_count[1][1] ),
    .Y(_0799_));
 sky130_fd_sc_hd__clkbuf_2 _1446_ (.A(\transfer_count[1][6] ),
    .X(_0800_));
 sky130_fd_sc_hd__nand2_1 _1447_ (.A(\transfer_count[1][7] ),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__nor4_2 _1448_ (.A(_0797_),
    .B(_0798_),
    .C(_0799_),
    .D(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__clkbuf_4 _1449_ (.A(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__and3_1 _1450_ (.A(\transfer_count[1][10] ),
    .B(\transfer_count[1][9] ),
    .C(\transfer_count[1][8] ),
    .X(_0804_));
 sky130_fd_sc_hd__and4_1 _1451_ (.A(\transfer_count[1][12] ),
    .B(\transfer_count[1][11] ),
    .C(_0803_),
    .D(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__xnor2_1 _1452_ (.A(\transfer_count[1][13] ),
    .B(_0805_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _1453_ (.A(\transfer_count[1][8] ),
    .B(_0803_),
    .Y(_0806_));
 sky130_fd_sc_hd__xor2_1 _1454_ (.A(\transfer_count[1][9] ),
    .B(_0806_),
    .X(_1051_));
 sky130_fd_sc_hd__and3_1 _1455_ (.A(\transfer_count[1][28] ),
    .B(\transfer_count[1][27] ),
    .C(\transfer_count[1][26] ),
    .X(_0807_));
 sky130_fd_sc_hd__inv_1 _1456_ (.A(\transfer_count[1][16] ),
    .Y(_0808_));
 sky130_fd_sc_hd__nand3_2 _1457_ (.A(\transfer_count[1][10] ),
    .B(\transfer_count[1][9] ),
    .C(\transfer_count[1][8] ),
    .Y(_0809_));
 sky130_fd_sc_hd__nand3_1 _1458_ (.A(\transfer_count[1][13] ),
    .B(\transfer_count[1][12] ),
    .C(\transfer_count[1][11] ),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(\transfer_count[1][14] ),
    .B(\transfer_count[1][15] ),
    .Y(_0811_));
 sky130_fd_sc_hd__nor4_4 _1460_ (.A(_0808_),
    .B(_0809_),
    .C(_0810_),
    .D(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_2 _1461_ (.A(\transfer_count[1][17] ),
    .X(_0813_));
 sky130_fd_sc_hd__nand4_1 _1462_ (.A(\transfer_count[1][20] ),
    .B(\transfer_count[1][19] ),
    .C(\transfer_count[1][18] ),
    .D(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(\transfer_count[1][22] ),
    .B(\transfer_count[1][21] ),
    .Y(_0815_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_0814_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__and2_0 _1465_ (.A(_0812_),
    .B(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__buf_4 _1466_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__and3_2 _1467_ (.A(\transfer_count[1][25] ),
    .B(\transfer_count[1][24] ),
    .C(\transfer_count[1][23] ),
    .X(_0819_));
 sky130_fd_sc_hd__nand4_4 _1468_ (.A(_0802_),
    .B(_0807_),
    .C(_0818_),
    .D(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__xor2_1 _1469_ (.A(\transfer_count[1][29] ),
    .B(_0820_),
    .X(_1063_));
 sky130_fd_sc_hd__inv_1 _1470_ (.A(\transfer_count[1][25] ),
    .Y(_0821_));
 sky130_fd_sc_hd__nand4_1 _1471_ (.A(\transfer_count[1][24] ),
    .B(\transfer_count[1][23] ),
    .C(_0803_),
    .D(_0818_),
    .Y(_0822_));
 sky130_fd_sc_hd__xnor2_1 _1472_ (.A(_0821_),
    .B(_0822_),
    .Y(_1075_));
 sky130_fd_sc_hd__nand2_2 _1473_ (.A(_0803_),
    .B(_0812_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(_0814_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__xnor2_1 _1475_ (.A(\transfer_count[1][21] ),
    .B(_0824_),
    .Y(_1087_));
 sky130_fd_sc_hd__xor2_1 _1476_ (.A(_0813_),
    .B(_0823_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_4 _1477_ (.A(\channel_state[1][0] ),
    .X(_0825_));
 sky130_fd_sc_hd__buf_2 _1478_ (.A(\channel_state[1][1] ),
    .X(_0826_));
 sky130_fd_sc_hd__nor2_2 _1479_ (.A(_0825_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand3_4 _1480_ (.A(net139),
    .B(\channel_state[1][2] ),
    .C(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__clkbuf_4 _1481_ (.A(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__a211oi_1 _1482_ (.A1(_1101_),
    .A2(_1103_),
    .B1(_1100_),
    .C1(_1097_),
    .Y(_0830_));
 sky130_fd_sc_hd__o21ai_0 _1483_ (.A1(_1098_),
    .A2(_1097_),
    .B1(_1095_),
    .Y(_0831_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(_1091_),
    .B(_1094_),
    .Y(_0832_));
 sky130_fd_sc_hd__o21a_1 _1485_ (.A1(_0830_),
    .A2(_0831_),
    .B1(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__o2111ai_1 _1486_ (.A1(_1092_),
    .A2(_1091_),
    .B1(_1083_),
    .C1(_1089_),
    .D1(_1086_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _1487_ (.A1(_1086_),
    .A2(_1088_),
    .B1(_1085_),
    .X(_0835_));
 sky130_fd_sc_hd__a21oi_1 _1488_ (.A1(_1083_),
    .A2(_0835_),
    .B1(_1082_),
    .Y(_0836_));
 sky130_fd_sc_hd__o21ai_1 _1489_ (.A1(_0833_),
    .A2(_0834_),
    .B1(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(_1059_),
    .B(_1062_),
    .Y(_0838_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_1065_),
    .B(_1068_),
    .Y(_0839_));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(_0838_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__a21oi_1 _1493_ (.A1(_1077_),
    .A2(_1079_),
    .B1(_1076_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_1071_),
    .B(_1074_),
    .Y(_0842_));
 sky130_fd_sc_hd__a21oi_1 _1495_ (.A1(_1071_),
    .A2(_1073_),
    .B1(_1070_),
    .Y(_0843_));
 sky130_fd_sc_hd__o21ai_2 _1496_ (.A1(_0841_),
    .A2(_0842_),
    .B1(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__a21oi_1 _1497_ (.A1(_1065_),
    .A2(_1067_),
    .B1(_1064_),
    .Y(_0845_));
 sky130_fd_sc_hd__a21oi_1 _1498_ (.A1(_1059_),
    .A2(_1061_),
    .B1(_1058_),
    .Y(_0846_));
 sky130_fd_sc_hd__o21ai_0 _1499_ (.A1(_0838_),
    .A2(_0845_),
    .B1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21oi_1 _1500_ (.A1(_0840_),
    .A2(_0844_),
    .B1(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__and3_1 _1501_ (.A(_1035_),
    .B(_1041_),
    .C(_1038_),
    .X(_0849_));
 sky130_fd_sc_hd__a211oi_1 _1502_ (.A1(_1053_),
    .A2(_1055_),
    .B1(_1052_),
    .C1(_1049_),
    .Y(_0850_));
 sky130_fd_sc_hd__o21ai_0 _1503_ (.A1(_1050_),
    .A2(_1049_),
    .B1(_1047_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(_1043_),
    .B(_1046_),
    .Y(_0852_));
 sky130_fd_sc_hd__o21ai_0 _1505_ (.A1(_0850_),
    .A2(_0851_),
    .B1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__o211ai_2 _1506_ (.A1(_1044_),
    .A2(_1043_),
    .B1(_0849_),
    .C1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2b_1 _1507_ (.A(_1410_),
    .B_N(_1416_),
    .Y(_0855_));
 sky130_fd_sc_hd__o211ai_1 _1508_ (.A1(_1415_),
    .A2(_0855_),
    .B1(_1419_),
    .C1(_1422_),
    .Y(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1509_ (.A1(_1419_),
    .A2(_1421_),
    .B1(_1418_),
    .Y(_0857_));
 sky130_fd_sc_hd__and4_1 _1510_ (.A(_1053_),
    .B(_1044_),
    .C(_1050_),
    .D(_1056_),
    .X(_0858_));
 sky130_fd_sc_hd__and4_1 _1511_ (.A(_1425_),
    .B(_1431_),
    .C(_1428_),
    .D(_1434_),
    .X(_0859_));
 sky130_fd_sc_hd__nand4_2 _1512_ (.A(_1047_),
    .B(_0858_),
    .C(_0849_),
    .D(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__a21o_1 _1513_ (.A1(_0856_),
    .A2(_0857_),
    .B1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__and3_1 _1514_ (.A(_1047_),
    .B(_0858_),
    .C(_0849_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_1 _1515_ (.A(_1425_),
    .B(_1428_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_1 _1516_ (.A1(_1431_),
    .A2(_1433_),
    .B1(_1430_),
    .Y(_0864_));
 sky130_fd_sc_hd__a21oi_1 _1517_ (.A1(_1425_),
    .A2(_1427_),
    .B1(_1424_),
    .Y(_0865_));
 sky130_fd_sc_hd__o21ai_1 _1518_ (.A1(_0863_),
    .A2(_0864_),
    .B1(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a21o_1 _1519_ (.A1(_1038_),
    .A2(_1040_),
    .B1(_1037_),
    .X(_0867_));
 sky130_fd_sc_hd__a221oi_1 _1520_ (.A1(_0862_),
    .A2(_0866_),
    .B1(_0867_),
    .B2(_1035_),
    .C1(_1034_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand4_1 _1521_ (.A(_0848_),
    .B(_0854_),
    .C(_0861_),
    .D(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand4_1 _1522_ (.A(_1083_),
    .B(_1089_),
    .C(_1101_),
    .D(_1086_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand4_1 _1523_ (.A(_1095_),
    .B(_1092_),
    .C(_1098_),
    .D(_1104_),
    .Y(_0871_));
 sky130_fd_sc_hd__nand4_1 _1524_ (.A(_1419_),
    .B(_1416_),
    .C(_1411_),
    .D(_1422_),
    .Y(_0872_));
 sky130_fd_sc_hd__nor4_1 _1525_ (.A(_0870_),
    .B(_0871_),
    .C(_0860_),
    .D(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _1526_ (.A(_1077_),
    .B(_1080_),
    .Y(_0874_));
 sky130_fd_sc_hd__nor2_1 _1527_ (.A(_0842_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _1528_ (.A(_0840_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__mux2i_1 _1529_ (.A0(_0873_),
    .A1(_0848_),
    .S(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__o21bai_1 _1530_ (.A1(_0870_),
    .A2(_0871_),
    .B1_N(_0847_),
    .Y(_0878_));
 sky130_fd_sc_hd__a211o_1 _1531_ (.A1(_0840_),
    .A2(_0844_),
    .B1(_0878_),
    .C1(_0837_),
    .X(_0879_));
 sky130_fd_sc_hd__o211a_1 _1532_ (.A1(_0837_),
    .A2(_0869_),
    .B1(_0877_),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__nor2b_1 _1533_ (.A(\channel_state[1][2] ),
    .B_N(net3),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_2 _1534_ (.A(net135),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nor3_1 _1535_ (.A(_0825_),
    .B(_0826_),
    .C(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__o22a_1 _1536_ (.A1(_0829_),
    .A2(_0880_),
    .B1(_0883_),
    .B2(net147),
    .X(_0005_));
 sky130_fd_sc_hd__buf_6 _1537_ (.A(\transfer_count[3][24] ),
    .X(_0884_));
 sky130_fd_sc_hd__and3_1 _1538_ (.A(\transfer_count[3][26] ),
    .B(\transfer_count[3][25] ),
    .C(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__nand3_1 _1539_ (.A(\transfer_count[3][28] ),
    .B(\transfer_count[3][27] ),
    .C(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__buf_6 _1540_ (.A(\transfer_count[3][23] ),
    .X(_0887_));
 sky130_fd_sc_hd__nand3_2 _1541_ (.A(\transfer_count[3][20] ),
    .B(\transfer_count[3][19] ),
    .C(\transfer_count[3][18] ),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _1542_ (.A(\transfer_count[3][22] ),
    .B(\transfer_count[3][21] ),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _1543_ (.A(_0888_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__nand4_4 _1544_ (.A(\transfer_count[3][5] ),
    .B(\transfer_count[3][4] ),
    .C(\transfer_count[3][3] ),
    .D(\transfer_count[3][2] ),
    .Y(_0891_));
 sky130_fd_sc_hd__nand3_1 _1545_ (.A(\transfer_count[3][6] ),
    .B(\transfer_count[3][1] ),
    .C(\transfer_count[3][0] ),
    .Y(_0892_));
 sky130_fd_sc_hd__nor2_2 _1546_ (.A(_0891_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__clkbuf_2 _1547_ (.A(\transfer_count[3][15] ),
    .X(_0894_));
 sky130_fd_sc_hd__nand3_2 _1548_ (.A(\transfer_count[3][17] ),
    .B(\transfer_count[3][16] ),
    .C(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand4_2 _1549_ (.A(\transfer_count[3][14] ),
    .B(\transfer_count[3][13] ),
    .C(\transfer_count[3][12] ),
    .D(\transfer_count[3][11] ),
    .Y(_0896_));
 sky130_fd_sc_hd__nand4_4 _1550_ (.A(\transfer_count[3][10] ),
    .B(\transfer_count[3][9] ),
    .C(\transfer_count[3][8] ),
    .D(\transfer_count[3][7] ),
    .Y(_0897_));
 sky130_fd_sc_hd__nor3_4 _1551_ (.A(_0895_),
    .B(_0896_),
    .C(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand4_2 _1552_ (.A(_0887_),
    .B(_0890_),
    .C(_0893_),
    .D(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__nor2_1 _1553_ (.A(_0886_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__xnor2_1 _1554_ (.A(\transfer_count[3][29] ),
    .B(_0900_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand3_1 _1555_ (.A(\transfer_count[3][26] ),
    .B(\transfer_count[3][25] ),
    .C(_0884_),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _1556_ (.A(_0901_),
    .B(_0899_),
    .Y(_0902_));
 sky130_fd_sc_hd__xnor2_1 _1557_ (.A(\transfer_count[3][27] ),
    .B(_0902_),
    .Y(_1117_));
 sky130_fd_sc_hd__or2_1 _1558_ (.A(_0895_),
    .B(_0896_),
    .X(_0903_));
 sky130_fd_sc_hd__or3_1 _1559_ (.A(_0897_),
    .B(_0891_),
    .C(_0892_),
    .X(_0904_));
 sky130_fd_sc_hd__buf_6 _1560_ (.A(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor4_4 _1561_ (.A(_0888_),
    .B(_0889_),
    .C(_0903_),
    .D(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__nand3_1 _1562_ (.A(_0884_),
    .B(_0887_),
    .C(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__xor2_1 _1563_ (.A(\transfer_count[3][25] ),
    .B(_0907_),
    .X(_1123_));
 sky130_fd_sc_hd__xnor2_1 _1564_ (.A(_0887_),
    .B(_0906_),
    .Y(_1129_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(_0888_),
    .B(_0895_),
    .Y(_0908_));
 sky130_fd_sc_hd__nor2_2 _1566_ (.A(_0896_),
    .B(_0905_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _1567_ (.A(_0908_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__xor2_1 _1568_ (.A(\transfer_count[3][21] ),
    .B(_0910_),
    .X(_1135_));
 sky130_fd_sc_hd__nor2_1 _1569_ (.A(_0903_),
    .B(_0905_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _1570_ (.A(\transfer_count[3][18] ),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__xor2_1 _1571_ (.A(\transfer_count[3][19] ),
    .B(_0912_),
    .X(_1141_));
 sky130_fd_sc_hd__xnor2_1 _1572_ (.A(_0894_),
    .B(_0909_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _1573_ (.A(\transfer_count[3][12] ),
    .B(\transfer_count[3][11] ),
    .Y(_0913_));
 sky130_fd_sc_hd__nor2_1 _1574_ (.A(_0913_),
    .B(_0905_),
    .Y(_0914_));
 sky130_fd_sc_hd__xnor2_1 _1575_ (.A(\transfer_count[3][13] ),
    .B(_0914_),
    .Y(_1159_));
 sky130_fd_sc_hd__inv_1 _1576_ (.A(\transfer_count[3][11] ),
    .Y(_0915_));
 sky130_fd_sc_hd__xnor2_1 _1577_ (.A(_0915_),
    .B(_0905_),
    .Y(_1165_));
 sky130_fd_sc_hd__and3_1 _1578_ (.A(\transfer_count[3][8] ),
    .B(\transfer_count[3][7] ),
    .C(_0893_),
    .X(_0916_));
 sky130_fd_sc_hd__xnor2_1 _1579_ (.A(\transfer_count[3][9] ),
    .B(_0916_),
    .Y(_1171_));
 sky130_fd_sc_hd__xnor2_1 _1580_ (.A(\transfer_count[3][7] ),
    .B(_0893_),
    .Y(_1177_));
 sky130_fd_sc_hd__and3_1 _1581_ (.A(\transfer_count[3][4] ),
    .B(\transfer_count[3][3] ),
    .C(\transfer_count[3][2] ),
    .X(_0917_));
 sky130_fd_sc_hd__nand3_1 _1582_ (.A(\transfer_count[3][1] ),
    .B(\transfer_count[3][0] ),
    .C(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__xor2_1 _1583_ (.A(\transfer_count[3][5] ),
    .B(_0918_),
    .X(_1183_));
 sky130_fd_sc_hd__nand3_1 _1584_ (.A(\transfer_count[3][2] ),
    .B(\transfer_count[3][1] ),
    .C(\transfer_count[3][0] ),
    .Y(_0919_));
 sky130_fd_sc_hd__xor2_1 _1585_ (.A(\transfer_count[3][3] ),
    .B(_0919_),
    .X(_1189_));
 sky130_fd_sc_hd__buf_2 _1586_ (.A(\channel_state[3][2] ),
    .X(_0920_));
 sky130_fd_sc_hd__nor2_1 _1587_ (.A(\channel_state[3][0] ),
    .B(\channel_state[3][1] ),
    .Y(_0921_));
 sky130_fd_sc_hd__nand3_2 _1588_ (.A(net141),
    .B(_0920_),
    .C(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__clkbuf_4 _1589_ (.A(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a21oi_1 _1590_ (.A1(_1115_),
    .A2(_1113_),
    .B1(_1112_),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_1 _1591_ (.A(_1107_),
    .B(_1110_),
    .Y(_0925_));
 sky130_fd_sc_hd__a21oi_1 _1592_ (.A1(_1107_),
    .A2(_1109_),
    .B1(_1106_),
    .Y(_0926_));
 sky130_fd_sc_hd__o21ai_0 _1593_ (.A1(_0924_),
    .A2(_0925_),
    .B1(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__nand4_1 _1594_ (.A(_1107_),
    .B(_1110_),
    .C(_1116_),
    .D(_1113_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand3_1 _1595_ (.A(_1127_),
    .B(_1122_),
    .C(_1125_),
    .Y(_0929_));
 sky130_fd_sc_hd__a21oi_1 _1596_ (.A1(_1122_),
    .A2(_1124_),
    .B1(_1121_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _1597_ (.A(_0929_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand4_1 _1598_ (.A(_1119_),
    .B(_1122_),
    .C(_1128_),
    .D(_1125_),
    .Y(_0932_));
 sky130_fd_sc_hd__a21oi_1 _1599_ (.A1(_1131_),
    .A2(_1133_),
    .B1(_1130_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_1 _1600_ (.A(_0932_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__a211oi_1 _1601_ (.A1(_1119_),
    .A2(_0931_),
    .B1(_0934_),
    .C1(_1118_),
    .Y(_0935_));
 sky130_fd_sc_hd__o21a_1 _1602_ (.A1(_1139_),
    .A2(_1140_),
    .B1(_1137_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2_1 _1603_ (.A(_1131_),
    .B(_1134_),
    .Y(_0937_));
 sky130_fd_sc_hd__nor3_1 _1604_ (.A(_0928_),
    .B(_0932_),
    .C(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a21oi_1 _1605_ (.A1(_1151_),
    .A2(_1149_),
    .B1(_1148_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _1606_ (.A(_1143_),
    .B(_1146_),
    .Y(_0940_));
 sky130_fd_sc_hd__a2111oi_0 _1607_ (.A1(_1143_),
    .A2(_1145_),
    .B1(_1136_),
    .C1(_1139_),
    .D1(_1142_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21ai_0 _1608_ (.A1(_0939_),
    .A2(_0940_),
    .B1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__o211ai_1 _1609_ (.A1(_1136_),
    .A2(_0936_),
    .B1(_0938_),
    .C1(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__o21ai_0 _1610_ (.A1(_0928_),
    .A2(_0935_),
    .B1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor3_1 _1611_ (.A(_0928_),
    .B(_0932_),
    .C(_0937_),
    .Y(_0945_));
 sky130_fd_sc_hd__and2_0 _1612_ (.A(_1143_),
    .B(_1140_),
    .X(_0946_));
 sky130_fd_sc_hd__and4_1 _1613_ (.A(_1146_),
    .B(_1149_),
    .C(_1152_),
    .D(_1137_),
    .X(_0947_));
 sky130_fd_sc_hd__nand4_1 _1614_ (.A(_1155_),
    .B(_1167_),
    .C(_1164_),
    .D(_1173_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand4_1 _1615_ (.A(_1158_),
    .B(_1170_),
    .C(_1176_),
    .D(_1161_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand4_1 _1616_ (.A(_1179_),
    .B(_1182_),
    .C(_1188_),
    .D(_1185_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand4_1 _1617_ (.A(_1191_),
    .B(_1199_),
    .C(_1203_),
    .D(_1194_),
    .Y(_0951_));
 sky130_fd_sc_hd__nor4_2 _1618_ (.A(_0948_),
    .B(_0949_),
    .C(_0950_),
    .D(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nand4_1 _1619_ (.A(_0945_),
    .B(_0946_),
    .C(_0947_),
    .D(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__o21a_1 _1620_ (.A1(_0927_),
    .A2(_0944_),
    .B1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2b_1 _1621_ (.A(_1202_),
    .B_N(_1199_),
    .Y(_0955_));
 sky130_fd_sc_hd__o211ai_1 _1622_ (.A1(_1198_),
    .A2(_0955_),
    .B1(_1191_),
    .C1(_1194_),
    .Y(_0956_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_1191_),
    .A2(_1193_),
    .B1(_1190_),
    .Y(_0957_));
 sky130_fd_sc_hd__a21oi_1 _1624_ (.A1(_0956_),
    .A2(_0957_),
    .B1(_0950_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand3_1 _1625_ (.A(_1187_),
    .B(_1182_),
    .C(_1185_),
    .Y(_0959_));
 sky130_fd_sc_hd__a21oi_1 _1626_ (.A1(_1182_),
    .A2(_1184_),
    .B1(_1181_),
    .Y(_0960_));
 sky130_fd_sc_hd__a21boi_0 _1627_ (.A1(_0959_),
    .A2(_0960_),
    .B1_N(_1179_),
    .Y(_0961_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0948_),
    .B(_0949_),
    .Y(_0962_));
 sky130_fd_sc_hd__o31ai_2 _1629_ (.A1(_1178_),
    .A2(_0958_),
    .A3(_0961_),
    .B1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a211oi_1 _1630_ (.A1(_1155_),
    .A2(_1157_),
    .B1(_1160_),
    .C1(_1163_),
    .Y(_0964_));
 sky130_fd_sc_hd__nand3_1 _1631_ (.A(_1175_),
    .B(_1170_),
    .C(_1173_),
    .Y(_0965_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(_1170_),
    .A2(_1172_),
    .B1(_1169_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(_1167_),
    .B(_1164_),
    .Y(_0967_));
 sky130_fd_sc_hd__a21o_1 _1634_ (.A1(_0965_),
    .A2(_0966_),
    .B1(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__nand2_1 _1635_ (.A(_1164_),
    .B(_1166_),
    .Y(_0969_));
 sky130_fd_sc_hd__o21a_1 _1636_ (.A1(_1161_),
    .A2(_1160_),
    .B1(_1158_),
    .X(_0970_));
 sky130_fd_sc_hd__o21ai_0 _1637_ (.A1(_1157_),
    .A2(_0970_),
    .B1(_1155_),
    .Y(_0971_));
 sky130_fd_sc_hd__a31oi_1 _1638_ (.A1(_0964_),
    .A2(_0968_),
    .A3(_0969_),
    .B1(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__nor2_1 _1639_ (.A(_1154_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand3_1 _1640_ (.A(_0945_),
    .B(_0946_),
    .C(_0947_),
    .Y(_0974_));
 sky130_fd_sc_hd__a211oi_4 _1641_ (.A1(_0963_),
    .A2(_0973_),
    .B1(_0952_),
    .C1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__buf_2 _1642_ (.A(\channel_state[3][0] ),
    .X(_0976_));
 sky130_fd_sc_hd__nor2b_1 _1643_ (.A(\channel_state[3][2] ),
    .B_N(net5),
    .Y(_0977_));
 sky130_fd_sc_hd__nand2_1 _1644_ (.A(net137),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__nor3_1 _1645_ (.A(_0976_),
    .B(\channel_state[3][1] ),
    .C(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__o32a_1 _1646_ (.A1(_0923_),
    .A2(_0954_),
    .A3(_0975_),
    .B1(_0979_),
    .B2(net149),
    .X(_0007_));
 sky130_fd_sc_hd__buf_2 _1647_ (.A(\channel_state[0][0] ),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_2 _1648_ (.A(\channel_state[0][1] ),
    .X(_0981_));
 sky130_fd_sc_hd__nor2b_1 _1649_ (.A(net134),
    .B_N(\channel_state[0][2] ),
    .Y(_0982_));
 sky130_fd_sc_hd__nand3b_1 _1650_ (.A_N(\channel_state[0][2] ),
    .B(net2),
    .C(net134),
    .Y(_0983_));
 sky130_fd_sc_hd__nor2_1 _1651_ (.A(_0981_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__a21oi_1 _1652_ (.A1(_0981_),
    .A2(_0982_),
    .B1(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__o21a_1 _1653_ (.A1(_0980_),
    .A2(_0985_),
    .B1(net154),
    .X(_0008_));
 sky130_fd_sc_hd__and3_1 _1654_ (.A(\transfer_count[0][2] ),
    .B(\transfer_count[0][1] ),
    .C(\transfer_count[0][0] ),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_2 _1655_ (.A(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__nand3_1 _1656_ (.A(\transfer_count[0][3] ),
    .B(\transfer_count[0][4] ),
    .C(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__xor2_1 _1657_ (.A(\transfer_count[0][5] ),
    .B(_0988_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_2 _1658_ (.A(\transfer_count[0][8] ),
    .X(_0989_));
 sky130_fd_sc_hd__nand3_1 _1659_ (.A(\transfer_count[0][10] ),
    .B(\transfer_count[0][9] ),
    .C(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__buf_2 _1660_ (.A(\transfer_count[0][7] ),
    .X(_0991_));
 sky130_fd_sc_hd__and3_2 _1661_ (.A(\transfer_count[0][3] ),
    .B(\transfer_count[0][5] ),
    .C(\transfer_count[0][4] ),
    .X(_0992_));
 sky130_fd_sc_hd__nand4_4 _1662_ (.A(\transfer_count[0][6] ),
    .B(_0991_),
    .C(_0987_),
    .D(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__nor2_1 _1663_ (.A(_0990_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand3_1 _1664_ (.A(\transfer_count[0][12] ),
    .B(\transfer_count[0][11] ),
    .C(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__xor2_1 _1665_ (.A(\transfer_count[0][13] ),
    .B(_0995_),
    .X(_1237_));
 sky130_fd_sc_hd__and3_1 _1666_ (.A(\transfer_count[0][6] ),
    .B(_0987_),
    .C(_0992_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_2 _1667_ (.A(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__nand3_1 _1668_ (.A(_0991_),
    .B(_0989_),
    .C(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__xor2_1 _1669_ (.A(\transfer_count[0][9] ),
    .B(_0998_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_2 _1670_ (.A(\transfer_count[0][22] ),
    .X(_0999_));
 sky130_fd_sc_hd__and4_1 _1671_ (.A(\transfer_count[0][25] ),
    .B(\transfer_count[0][24] ),
    .C(\transfer_count[0][23] ),
    .D(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1672_ (.A(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__and4_1 _1673_ (.A(\transfer_count[0][28] ),
    .B(\transfer_count[0][27] ),
    .C(\transfer_count[0][26] ),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__buf_2 _1674_ (.A(\transfer_count[0][16] ),
    .X(_1003_));
 sky130_fd_sc_hd__and3_1 _1675_ (.A(\transfer_count[0][18] ),
    .B(\transfer_count[0][17] ),
    .C(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__nand4_4 _1676_ (.A(\transfer_count[0][21] ),
    .B(\transfer_count[0][20] ),
    .C(\transfer_count[0][19] ),
    .D(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__and3_2 _1677_ (.A(\transfer_count[0][10] ),
    .B(\transfer_count[0][9] ),
    .C(_0989_),
    .X(_1006_));
 sky130_fd_sc_hd__and3_1 _1678_ (.A(\transfer_count[0][13] ),
    .B(\transfer_count[0][12] ),
    .C(\transfer_count[0][11] ),
    .X(_1007_));
 sky130_fd_sc_hd__nand4_4 _1679_ (.A(\transfer_count[0][14] ),
    .B(\transfer_count[0][15] ),
    .C(_1006_),
    .D(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__nor3_4 _1680_ (.A(_0993_),
    .B(_1005_),
    .C(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2_1 _1681_ (.A(_1002_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__xor2_1 _1682_ (.A(\transfer_count[0][29] ),
    .B(_1010_),
    .X(_1261_));
 sky130_fd_sc_hd__and3_1 _1683_ (.A(\transfer_count[0][24] ),
    .B(\transfer_count[0][23] ),
    .C(_0999_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(_1011_),
    .B(_1009_),
    .Y(_1012_));
 sky130_fd_sc_hd__xor2_1 _1685_ (.A(\transfer_count[0][25] ),
    .B(_1012_),
    .X(_1273_));
 sky130_fd_sc_hd__and3_1 _1686_ (.A(\transfer_count[0][20] ),
    .B(\transfer_count[0][19] ),
    .C(_1004_),
    .X(_1013_));
 sky130_fd_sc_hd__nand3_1 _1687_ (.A(\transfer_count[0][14] ),
    .B(_1006_),
    .C(_1007_),
    .Y(_1014_));
 sky130_fd_sc_hd__nor2_2 _1688_ (.A(_0993_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__and3_1 _1689_ (.A(\transfer_count[0][15] ),
    .B(_1013_),
    .C(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__xnor2_1 _1690_ (.A(\transfer_count[0][21] ),
    .B(_1016_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand3_1 _1691_ (.A(\transfer_count[0][15] ),
    .B(_1003_),
    .C(_1015_),
    .Y(_0146_));
 sky130_fd_sc_hd__xor2_1 _1692_ (.A(\transfer_count[0][17] ),
    .B(_0146_),
    .X(_1297_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(net138),
    .B(\channel_state[0][2] ),
    .Y(_0147_));
 sky130_fd_sc_hd__nor3_1 _1694_ (.A(_0980_),
    .B(_0981_),
    .C(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__clkbuf_4 _1695_ (.A(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_4 _1696_ (.A(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__nand4_2 _1697_ (.A(_1257_),
    .B(_1263_),
    .C(_1260_),
    .D(_1266_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand4_1 _1698_ (.A(_1269_),
    .B(_1275_),
    .C(_1272_),
    .D(_1278_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand3_1 _1699_ (.A(_1281_),
    .B(_1287_),
    .C(_1284_),
    .Y(_0153_));
 sky130_fd_sc_hd__nor3_2 _1700_ (.A(_0151_),
    .B(_0152_),
    .C(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__and3_1 _1701_ (.A(_1293_),
    .B(_1290_),
    .C(_1296_),
    .X(_0155_));
 sky130_fd_sc_hd__nand4_2 _1702_ (.A(_1299_),
    .B(_1302_),
    .C(_0154_),
    .D(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand3_1 _1703_ (.A(_1233_),
    .B(_1239_),
    .C(_1236_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand4_1 _1704_ (.A(_1251_),
    .B(_1242_),
    .C(_1248_),
    .D(_1254_),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2_1 _1705_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand3_1 _1706_ (.A(_1215_),
    .B(_1218_),
    .C(_1230_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand4_1 _1707_ (.A(_1207_),
    .B(_1221_),
    .C(_1227_),
    .D(_1224_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _1708_ (.A(_0160_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand4_2 _1709_ (.A(_1212_),
    .B(_1245_),
    .C(_0159_),
    .D(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__a21o_1 _1710_ (.A1(_1293_),
    .A2(_1295_),
    .B1(_1292_),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_1 _1711_ (.A1(_1299_),
    .A2(_1301_),
    .B1(_1298_),
    .X(_0165_));
 sky130_fd_sc_hd__a221oi_1 _1712_ (.A1(_1290_),
    .A2(_0164_),
    .B1(_0165_),
    .B2(_0155_),
    .C1(_1289_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2b_1 _1713_ (.A(_0166_),
    .B_N(_0154_),
    .Y(_0167_));
 sky130_fd_sc_hd__a21o_1 _1714_ (.A1(_1275_),
    .A2(_1277_),
    .B1(_1274_),
    .X(_0168_));
 sky130_fd_sc_hd__nand3_1 _1715_ (.A(_1269_),
    .B(_1272_),
    .C(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__a21oi_1 _1716_ (.A1(_1269_),
    .A2(_1271_),
    .B1(_1268_),
    .Y(_0170_));
 sky130_fd_sc_hd__a21oi_1 _1717_ (.A1(_0169_),
    .A2(_0170_),
    .B1(_0151_),
    .Y(_0171_));
 sky130_fd_sc_hd__a21o_1 _1718_ (.A1(_1284_),
    .A2(_1286_),
    .B1(_1283_),
    .X(_0172_));
 sky130_fd_sc_hd__a21oi_1 _1719_ (.A1(_1281_),
    .A2(_0172_),
    .B1(_1280_),
    .Y(_0173_));
 sky130_fd_sc_hd__a211oi_1 _1720_ (.A1(_1263_),
    .A2(_1265_),
    .B1(_1262_),
    .C1(_1259_),
    .Y(_0174_));
 sky130_fd_sc_hd__o21ai_0 _1721_ (.A1(_1260_),
    .A2(_1259_),
    .B1(_1257_),
    .Y(_0175_));
 sky130_fd_sc_hd__o32ai_1 _1722_ (.A1(_0151_),
    .A2(_0152_),
    .A3(_0173_),
    .B1(_0174_),
    .B2(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__or4_2 _1723_ (.A(_1256_),
    .B(_0167_),
    .C(_0171_),
    .D(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_1 _1724_ (.A1(_1236_),
    .A2(_1238_),
    .B1(_1235_),
    .X(_0178_));
 sky130_fd_sc_hd__a21oi_1 _1725_ (.A1(_1233_),
    .A2(_0178_),
    .B1(_1232_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21o_1 _1726_ (.A1(_1224_),
    .A2(_1226_),
    .B1(_1223_),
    .X(_0180_));
 sky130_fd_sc_hd__a211o_1 _1727_ (.A1(_1221_),
    .A2(_0180_),
    .B1(_1229_),
    .C1(_1220_),
    .X(_0181_));
 sky130_fd_sc_hd__inv_1 _1728_ (.A(_1211_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2b_1 _1729_ (.A_N(_1206_),
    .B(_1212_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _1730_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_0160_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _1731_ (.A1(_1215_),
    .A2(_1217_),
    .B1(_1214_),
    .Y(_0185_));
 sky130_fd_sc_hd__nor2b_1 _1732_ (.A(_0185_),
    .B_N(_1230_),
    .Y(_0186_));
 sky130_fd_sc_hd__nor3_1 _1733_ (.A(_1227_),
    .B(_1223_),
    .C(_1226_),
    .Y(_0187_));
 sky130_fd_sc_hd__o21ai_0 _1734_ (.A1(_1224_),
    .A2(_1223_),
    .B1(_1221_),
    .Y(_0188_));
 sky130_fd_sc_hd__o21bai_1 _1735_ (.A1(_0187_),
    .A2(_0188_),
    .B1_N(_1220_),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_1245_),
    .B(_1254_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand3_1 _1737_ (.A(_1251_),
    .B(_1242_),
    .C(_1248_),
    .Y(_0191_));
 sky130_fd_sc_hd__nor3_1 _1738_ (.A(_0157_),
    .B(_0190_),
    .C(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__o311ai_2 _1739_ (.A1(_0181_),
    .A2(_0184_),
    .A3(_0186_),
    .B1(_0189_),
    .C1(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__a211oi_1 _1740_ (.A1(_1251_),
    .A2(_1253_),
    .B1(_1250_),
    .C1(_1247_),
    .Y(_0194_));
 sky130_fd_sc_hd__o21ai_0 _1741_ (.A1(_1248_),
    .A2(_1247_),
    .B1(_1245_),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_1 _1742_ (.A(_0194_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _1743_ (.A(_1242_),
    .B(_1241_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _1744_ (.A(_0157_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__o31ai_1 _1745_ (.A1(_1241_),
    .A2(_1244_),
    .A3(_0196_),
    .B1(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__a31oi_2 _1746_ (.A1(_0179_),
    .A2(_0193_),
    .A3(_0199_),
    .B1(_0156_),
    .Y(_0200_));
 sky130_fd_sc_hd__o22ai_4 _1747_ (.A1(_0156_),
    .A2(_0163_),
    .B1(_0177_),
    .B2(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor3_2 _1748_ (.A(_0980_),
    .B(_0981_),
    .C(_0983_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_1 _1749_ (.A(net146),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_1 _1750_ (.A1(_0150_),
    .A2(_0201_),
    .B1(_0203_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_1 _1751_ (.A(\transfer_count[3][0] ),
    .Y(_1201_));
 sky130_fd_sc_hd__clkbuf_4 _1752_ (.A(_0923_),
    .X(_0204_));
 sky130_fd_sc_hd__and3_1 _1753_ (.A(net141),
    .B(\channel_state[3][2] ),
    .C(_0921_),
    .X(_0205_));
 sky130_fd_sc_hd__buf_2 _1754_ (.A(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _1755_ (.A(_0206_),
    .B(_0979_),
    .Y(_0207_));
 sky130_fd_sc_hd__clkbuf_4 _1756_ (.A(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _1757_ (.A(\transfer_count[3][0] ),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__o21ai_0 _1758_ (.A1(\transfer_count[3][0] ),
    .A2(_0204_),
    .B1(_0209_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_1 _1759_ (.A(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _1760_ (.A(\transfer_count[3][1] ),
    .B(_0208_),
    .Y(_0210_));
 sky130_fd_sc_hd__o21ai_0 _1761_ (.A1(_1197_),
    .A2(_0204_),
    .B1(_0210_),
    .Y(_0120_));
 sky130_fd_sc_hd__clkbuf_2 _1762_ (.A(_1195_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_4 _1763_ (.A(_0206_),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(_0211_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__clkbuf_4 _1765_ (.A(_0922_),
    .X(_0214_));
 sky130_fd_sc_hd__o31ai_2 _1766_ (.A1(_0976_),
    .A2(\channel_state[3][1] ),
    .A3(_0978_),
    .B1(_0922_),
    .Y(_0215_));
 sky130_fd_sc_hd__clkbuf_4 _1767_ (.A(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ai_0 _1768_ (.A1(_0211_),
    .A2(_0214_),
    .B1(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1769_ (.A(\transfer_count[3][2] ),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__o21ai_0 _1770_ (.A1(\transfer_count[3][2] ),
    .A2(_0213_),
    .B1(_0218_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(\transfer_count[3][3] ),
    .B(_0208_),
    .Y(_0219_));
 sky130_fd_sc_hd__o21ai_0 _1772_ (.A1(_1189_),
    .A2(_0204_),
    .B1(_0219_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand3_1 _1773_ (.A(\transfer_count[3][3] ),
    .B(\transfer_count[3][2] ),
    .C(_0211_),
    .Y(_0220_));
 sky130_fd_sc_hd__xor2_1 _1774_ (.A(\transfer_count[3][4] ),
    .B(_0220_),
    .X(_1186_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(\transfer_count[3][4] ),
    .B(_0208_),
    .Y(_0221_));
 sky130_fd_sc_hd__o21ai_0 _1776_ (.A1(_0204_),
    .A2(_1186_),
    .B1(_0221_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _1777_ (.A(\transfer_count[3][5] ),
    .B(_0208_),
    .Y(_0222_));
 sky130_fd_sc_hd__o21ai_0 _1778_ (.A1(_1183_),
    .A2(_0204_),
    .B1(_0222_),
    .Y(_0136_));
 sky130_fd_sc_hd__clkbuf_4 _1779_ (.A(_0923_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_0 _1780_ (.A(\transfer_count[3][5] ),
    .B(_0917_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _1781_ (.A(_0211_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__buf_4 _1782_ (.A(_0207_),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_1 _1783_ (.A1(_0211_),
    .A2(_0224_),
    .B1(_0214_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_0 _1784_ (.A1(_0226_),
    .A2(_0227_),
    .B1(\transfer_count[3][6] ),
    .Y(_0228_));
 sky130_fd_sc_hd__o31ai_1 _1785_ (.A1(\transfer_count[3][6] ),
    .A2(_0223_),
    .A3(_0225_),
    .B1(_0228_),
    .Y(_0137_));
 sky130_fd_sc_hd__nor2_1 _1786_ (.A(_0893_),
    .B(_0214_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_0 _1787_ (.A1(_0226_),
    .A2(_0229_),
    .B1(\transfer_count[3][7] ),
    .Y(_0230_));
 sky130_fd_sc_hd__o41ai_1 _1788_ (.A1(\transfer_count[3][7] ),
    .A2(_0891_),
    .A3(_0892_),
    .A4(_0223_),
    .B1(_0230_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _1789_ (.A(\transfer_count[3][6] ),
    .B(_0211_),
    .Y(_0231_));
 sky130_fd_sc_hd__nor2_2 _1790_ (.A(_0891_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(\transfer_count[3][7] ),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__xor2_1 _1792_ (.A(\transfer_count[3][8] ),
    .B(_0233_),
    .X(_1174_));
 sky130_fd_sc_hd__nand2_1 _1793_ (.A(\transfer_count[3][8] ),
    .B(_0208_),
    .Y(_0234_));
 sky130_fd_sc_hd__o21ai_0 _1794_ (.A1(_0204_),
    .A2(_1174_),
    .B1(_0234_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _1795_ (.A(\transfer_count[3][9] ),
    .B(_0208_),
    .Y(_0235_));
 sky130_fd_sc_hd__o21ai_0 _1796_ (.A1(_1171_),
    .A2(_0204_),
    .B1(_0235_),
    .Y(_0140_));
 sky130_fd_sc_hd__and4_1 _1797_ (.A(\transfer_count[3][9] ),
    .B(\transfer_count[3][8] ),
    .C(\transfer_count[3][7] ),
    .D(_0232_),
    .X(_0236_));
 sky130_fd_sc_hd__xnor2_1 _1798_ (.A(\transfer_count[3][10] ),
    .B(_0236_),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_1 _1799_ (.A(\transfer_count[3][10] ),
    .B(_0208_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_0 _1800_ (.A1(_0204_),
    .A2(_1168_),
    .B1(_0237_),
    .Y(_0110_));
 sky130_fd_sc_hd__a21oi_1 _1801_ (.A1(_0905_),
    .A2(_0206_),
    .B1(_0207_),
    .Y(_0238_));
 sky130_fd_sc_hd__or3_1 _1802_ (.A(\transfer_count[3][11] ),
    .B(_0905_),
    .C(_0922_),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_0 _1803_ (.A1(_0915_),
    .A2(_0238_),
    .B1(_0239_),
    .Y(_0111_));
 sky130_fd_sc_hd__nor4_1 _1804_ (.A(_0915_),
    .B(_0897_),
    .C(_0891_),
    .D(_0231_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_1 _1805_ (.A(\transfer_count[3][12] ),
    .B(_0240_),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_1 _1806_ (.A(\transfer_count[3][12] ),
    .B(_0208_),
    .Y(_0241_));
 sky130_fd_sc_hd__o21ai_0 _1807_ (.A1(_0204_),
    .A2(_1162_),
    .B1(_0241_),
    .Y(_0112_));
 sky130_fd_sc_hd__nand2_1 _1808_ (.A(_0914_),
    .B(_0212_),
    .Y(_0242_));
 sky130_fd_sc_hd__o21ai_0 _1809_ (.A1(_0914_),
    .A2(_0214_),
    .B1(_0216_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _1810_ (.A(\transfer_count[3][13] ),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__o21ai_0 _1811_ (.A1(\transfer_count[3][13] ),
    .A2(_0242_),
    .B1(_0244_),
    .Y(_0113_));
 sky130_fd_sc_hd__nand3_1 _1812_ (.A(\transfer_count[3][13] ),
    .B(\transfer_count[3][12] ),
    .C(\transfer_count[3][11] ),
    .Y(_0245_));
 sky130_fd_sc_hd__nor4_2 _1813_ (.A(_0245_),
    .B(_0897_),
    .C(_0891_),
    .D(_0231_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand2_1 _1814_ (.A(_0212_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__o21ai_0 _1815_ (.A1(_0923_),
    .A2(_0246_),
    .B1(_0216_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _1816_ (.A(\transfer_count[3][14] ),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__o21ai_0 _1817_ (.A1(\transfer_count[3][14] ),
    .A2(_0247_),
    .B1(_0249_),
    .Y(_0114_));
 sky130_fd_sc_hd__o21ai_0 _1818_ (.A1(_0909_),
    .A2(_0923_),
    .B1(_0215_),
    .Y(_0250_));
 sky130_fd_sc_hd__nor2_1 _1819_ (.A(_0894_),
    .B(_0214_),
    .Y(_0251_));
 sky130_fd_sc_hd__a22o_1 _1820_ (.A1(_0894_),
    .A2(_0250_),
    .B1(_0251_),
    .B2(_0909_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _1821_ (.A(_0894_),
    .B(\transfer_count[3][14] ),
    .C(_0246_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _1822_ (.A(_0212_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__o21ai_0 _1823_ (.A1(_0923_),
    .A2(_0252_),
    .B1(_0216_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _1824_ (.A(\transfer_count[3][16] ),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__o21ai_0 _1825_ (.A1(\transfer_count[3][16] ),
    .A2(_0253_),
    .B1(_0255_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand3_1 _1826_ (.A(\transfer_count[3][16] ),
    .B(_0894_),
    .C(_0909_),
    .Y(_0256_));
 sky130_fd_sc_hd__a31oi_1 _1827_ (.A1(\transfer_count[3][16] ),
    .A2(_0894_),
    .A3(_0909_),
    .B1(_0923_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21ai_0 _1828_ (.A1(_0226_),
    .A2(_0257_),
    .B1(\transfer_count[3][17] ),
    .Y(_0258_));
 sky130_fd_sc_hd__o31ai_1 _1829_ (.A1(\transfer_count[3][17] ),
    .A2(_0223_),
    .A3(_0256_),
    .B1(_0258_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _1830_ (.A(_0898_),
    .B(_0232_),
    .Y(_0259_));
 sky130_fd_sc_hd__a21oi_1 _1831_ (.A1(_0898_),
    .A2(_0232_),
    .B1(_0214_),
    .Y(_0260_));
 sky130_fd_sc_hd__o21ai_0 _1832_ (.A1(_0226_),
    .A2(_0260_),
    .B1(\transfer_count[3][18] ),
    .Y(_0261_));
 sky130_fd_sc_hd__o31ai_1 _1833_ (.A1(\transfer_count[3][18] ),
    .A2(_0223_),
    .A3(_0259_),
    .B1(_0261_),
    .Y(_0118_));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(\transfer_count[3][19] ),
    .B(_0226_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_0 _1835_ (.A1(_1141_),
    .A2(_0204_),
    .B1(_0262_),
    .Y(_0119_));
 sky130_fd_sc_hd__and4_1 _1836_ (.A(\transfer_count[3][19] ),
    .B(\transfer_count[3][18] ),
    .C(_0898_),
    .D(_0232_),
    .X(_0263_));
 sky130_fd_sc_hd__o21ai_0 _1837_ (.A1(_0923_),
    .A2(_0263_),
    .B1(_0215_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(\transfer_count[3][20] ),
    .B(_0214_),
    .Y(_0265_));
 sky130_fd_sc_hd__a22o_1 _1839_ (.A1(\transfer_count[3][20] ),
    .A2(_0264_),
    .B1(_0265_),
    .B2(_0263_),
    .X(_0121_));
 sky130_fd_sc_hd__a21oi_1 _1840_ (.A1(_0908_),
    .A2(_0909_),
    .B1(_0214_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_0 _1841_ (.A1(_0226_),
    .A2(_0266_),
    .B1(\transfer_count[3][21] ),
    .Y(_0267_));
 sky130_fd_sc_hd__o31ai_1 _1842_ (.A1(\transfer_count[3][21] ),
    .A2(_0910_),
    .A3(_0223_),
    .B1(_0267_),
    .Y(_0122_));
 sky130_fd_sc_hd__and3_1 _1843_ (.A(\transfer_count[3][21] ),
    .B(\transfer_count[3][20] ),
    .C(_0263_),
    .X(_0268_));
 sky130_fd_sc_hd__nand2b_1 _1844_ (.A_N(_0268_),
    .B(_0206_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21oi_1 _1845_ (.A1(_0212_),
    .A2(_0268_),
    .B1(\transfer_count[3][22] ),
    .Y(_0270_));
 sky130_fd_sc_hd__a31oi_1 _1846_ (.A1(\transfer_count[3][22] ),
    .A2(_0216_),
    .A3(_0269_),
    .B1(_0270_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _1847_ (.A(_0906_),
    .B(_0212_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21ai_0 _1848_ (.A1(_0906_),
    .A2(_0214_),
    .B1(_0216_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _1849_ (.A(_0887_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ai_0 _1850_ (.A1(_0887_),
    .A2(_0271_),
    .B1(_0273_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand4_4 _1851_ (.A(_0887_),
    .B(_0890_),
    .C(_0898_),
    .D(_0232_),
    .Y(_0274_));
 sky130_fd_sc_hd__and2_0 _1852_ (.A(_0206_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__o21ai_0 _1853_ (.A1(_0226_),
    .A2(_0275_),
    .B1(_0884_),
    .Y(_0276_));
 sky130_fd_sc_hd__o31ai_1 _1854_ (.A1(_0884_),
    .A2(_0223_),
    .A3(_0274_),
    .B1(_0276_),
    .Y(_0125_));
 sky130_fd_sc_hd__a31oi_1 _1855_ (.A1(_0884_),
    .A2(_0887_),
    .A3(_0906_),
    .B1(_0923_),
    .Y(_0277_));
 sky130_fd_sc_hd__o21ai_0 _1856_ (.A1(_0226_),
    .A2(_0277_),
    .B1(\transfer_count[3][25] ),
    .Y(_0278_));
 sky130_fd_sc_hd__o31ai_1 _1857_ (.A1(\transfer_count[3][25] ),
    .A2(_0907_),
    .A3(_0223_),
    .B1(_0278_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _1858_ (.A(\transfer_count[3][25] ),
    .B(_0884_),
    .Y(_0279_));
 sky130_fd_sc_hd__o21ai_0 _1859_ (.A1(_0279_),
    .A2(_0274_),
    .B1(_0206_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _1860_ (.A(_0279_),
    .B(_0274_),
    .Y(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1861_ (.A1(_0212_),
    .A2(_0281_),
    .B1(\transfer_count[3][26] ),
    .Y(_0282_));
 sky130_fd_sc_hd__a31oi_1 _1862_ (.A1(\transfer_count[3][26] ),
    .A2(_0216_),
    .A3(_0280_),
    .B1(_0282_),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _1863_ (.A(_0887_),
    .B(_0906_),
    .Y(_0283_));
 sky130_fd_sc_hd__a31oi_1 _1864_ (.A1(_0887_),
    .A2(_0885_),
    .A3(_0906_),
    .B1(_0214_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_0 _1865_ (.A1(_0226_),
    .A2(_0284_),
    .B1(\transfer_count[3][27] ),
    .Y(_0285_));
 sky130_fd_sc_hd__o41ai_1 _1866_ (.A1(\transfer_count[3][27] ),
    .A2(_0901_),
    .A3(_0283_),
    .A4(_0223_),
    .B1(_0285_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(\transfer_count[3][27] ),
    .B(_0885_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_0 _1868_ (.A1(_0286_),
    .A2(_0274_),
    .B1(_0206_),
    .Y(_0287_));
 sky130_fd_sc_hd__nor2_1 _1869_ (.A(_0286_),
    .B(_0274_),
    .Y(_0288_));
 sky130_fd_sc_hd__a21oi_1 _1870_ (.A1(_0212_),
    .A2(_0288_),
    .B1(\transfer_count[3][28] ),
    .Y(_0289_));
 sky130_fd_sc_hd__a31oi_1 _1871_ (.A1(\transfer_count[3][28] ),
    .A2(_0216_),
    .A3(_0287_),
    .B1(_0289_),
    .Y(_0129_));
 sky130_fd_sc_hd__and3_1 _1872_ (.A(\transfer_count[3][28] ),
    .B(\transfer_count[3][27] ),
    .C(_0885_),
    .X(_0290_));
 sky130_fd_sc_hd__a31oi_1 _1873_ (.A1(_0887_),
    .A2(_0290_),
    .A3(_0906_),
    .B1(_0923_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21ai_0 _1874_ (.A1(_0226_),
    .A2(_0291_),
    .B1(\transfer_count[3][29] ),
    .Y(_0292_));
 sky130_fd_sc_hd__o41ai_1 _1875_ (.A1(\transfer_count[3][29] ),
    .A2(_0886_),
    .A3(_0283_),
    .A4(_0223_),
    .B1(_0292_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _1876_ (.A(\transfer_count[3][29] ),
    .B(_0290_),
    .Y(_0293_));
 sky130_fd_sc_hd__o21ai_0 _1877_ (.A1(_0274_),
    .A2(_0293_),
    .B1(_0206_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _1878_ (.A(_0274_),
    .B(_0293_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1879_ (.A1(_0212_),
    .A2(_0295_),
    .B1(\transfer_count[3][30] ),
    .Y(_0296_));
 sky130_fd_sc_hd__a31oi_1 _1880_ (.A1(\transfer_count[3][30] ),
    .A2(_0216_),
    .A3(_0294_),
    .B1(_0296_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand3_1 _1881_ (.A(\transfer_count[3][30] ),
    .B(\transfer_count[3][29] ),
    .C(_0290_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_0 _1882_ (.A1(_0899_),
    .A2(_0297_),
    .B1(_0206_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(_0899_),
    .B(_0297_),
    .Y(_0299_));
 sky130_fd_sc_hd__a21oi_1 _1884_ (.A1(_0212_),
    .A2(_0299_),
    .B1(\transfer_count[3][31] ),
    .Y(_0300_));
 sky130_fd_sc_hd__a31oi_1 _1885_ (.A1(\transfer_count[3][31] ),
    .A2(_0216_),
    .A3(_0298_),
    .B1(_0300_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_1 _1886_ (.A(\transfer_count[2][0] ),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2b_1 _1887_ (.A_N(\channel_state[2][0] ),
    .B(\channel_state[2][2] ),
    .Y(_0301_));
 sky130_fd_sc_hd__nor2_1 _1888_ (.A(\channel_state[2][1] ),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_2 _1889_ (.A(net140),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__buf_2 _1890_ (.A(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__and2_0 _1891_ (.A(net140),
    .B(_0302_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_2 _1892_ (.A(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__inv_1 _1893_ (.A(\channel_state[2][0] ),
    .Y(_0307_));
 sky130_fd_sc_hd__buf_2 _1894_ (.A(\channel_state[2][2] ),
    .X(_0308_));
 sky130_fd_sc_hd__nor2b_1 _1895_ (.A(_0308_),
    .B_N(net4),
    .Y(_0309_));
 sky130_fd_sc_hd__and3_1 _1896_ (.A(_0307_),
    .B(net136),
    .C(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__nor2b_1 _1897_ (.A(\channel_state[2][1] ),
    .B_N(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_2 _1898_ (.A(_0306_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__buf_2 _1899_ (.A(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _1900_ (.A(\transfer_count[2][0] ),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__o21ai_0 _1901_ (.A1(\transfer_count[2][0] ),
    .A2(_0304_),
    .B1(_0314_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _1902_ (.A(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__nand2_1 _1903_ (.A(\transfer_count[2][1] ),
    .B(_0313_),
    .Y(_0315_));
 sky130_fd_sc_hd__o21ai_0 _1904_ (.A1(_1401_),
    .A2(_0304_),
    .B1(_0315_),
    .Y(_0088_));
 sky130_fd_sc_hd__clkbuf_4 _1905_ (.A(_0306_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _1906_ (.A(_1399_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__clkbuf_4 _1907_ (.A(_0312_),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_4 _1908_ (.A(_0303_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _1909_ (.A(_1399_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_0 _1910_ (.A1(_0318_),
    .A2(_0320_),
    .B1(\transfer_count[2][2] ),
    .Y(_0321_));
 sky130_fd_sc_hd__o21ai_0 _1911_ (.A1(\transfer_count[2][2] ),
    .A2(_0317_),
    .B1(_0321_),
    .Y(_0099_));
 sky130_fd_sc_hd__nand3_1 _1912_ (.A(\transfer_count[2][0] ),
    .B(\transfer_count[2][1] ),
    .C(\transfer_count[2][2] ),
    .Y(_0322_));
 sky130_fd_sc_hd__xor2_1 _1913_ (.A(\transfer_count[2][3] ),
    .B(_0322_),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_1 _1914_ (.A(\transfer_count[2][3] ),
    .B(_0313_),
    .Y(_0323_));
 sky130_fd_sc_hd__o21ai_0 _1915_ (.A1(_0304_),
    .A2(_1393_),
    .B1(_0323_),
    .Y(_0102_));
 sky130_fd_sc_hd__buf_4 _1916_ (.A(\transfer_count[2][4] ),
    .X(_0324_));
 sky130_fd_sc_hd__and3_1 _1917_ (.A(\transfer_count[2][2] ),
    .B(\transfer_count[2][3] ),
    .C(_1399_),
    .X(_0325_));
 sky130_fd_sc_hd__xnor2_2 _1918_ (.A(_0324_),
    .B(_0325_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(_0324_),
    .B(_0313_),
    .Y(_0326_));
 sky130_fd_sc_hd__o21ai_0 _1920_ (.A1(_0304_),
    .A2(_1390_),
    .B1(_0326_),
    .Y(_0103_));
 sky130_fd_sc_hd__and4_1 _1921_ (.A(\transfer_count[2][0] ),
    .B(\transfer_count[2][1] ),
    .C(\transfer_count[2][2] ),
    .D(\transfer_count[2][3] ),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(_0324_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _1923_ (.A(\transfer_count[2][5] ),
    .B(_0328_),
    .X(_1387_));
 sky130_fd_sc_hd__a21oi_1 _1924_ (.A1(_0324_),
    .A2(_0327_),
    .B1(_0319_),
    .Y(_0329_));
 sky130_fd_sc_hd__o21ai_0 _1925_ (.A1(_0313_),
    .A2(_0329_),
    .B1(\transfer_count[2][5] ),
    .Y(_0330_));
 sky130_fd_sc_hd__o31ai_1 _1926_ (.A1(\transfer_count[2][5] ),
    .A2(_0304_),
    .A3(_0328_),
    .B1(_0330_),
    .Y(_0104_));
 sky130_fd_sc_hd__and3_1 _1927_ (.A(_0324_),
    .B(\transfer_count[2][5] ),
    .C(_0325_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(_0316_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(_0319_),
    .B(_0331_),
    .Y(_0333_));
 sky130_fd_sc_hd__o21ai_0 _1930_ (.A1(_0318_),
    .A2(_0333_),
    .B1(\transfer_count[2][6] ),
    .Y(_0334_));
 sky130_fd_sc_hd__o21ai_0 _1931_ (.A1(\transfer_count[2][6] ),
    .A2(_0332_),
    .B1(_0334_),
    .Y(_0105_));
 sky130_fd_sc_hd__and2_1 _1932_ (.A(\transfer_count[2][5] ),
    .B(\transfer_count[2][6] ),
    .X(_0335_));
 sky130_fd_sc_hd__and3_1 _1933_ (.A(_0324_),
    .B(_0327_),
    .C(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1934_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__xnor2_1 _1935_ (.A(\transfer_count[2][7] ),
    .B(_0337_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand3_2 _1936_ (.A(_0324_),
    .B(_0327_),
    .C(_0335_),
    .Y(_0338_));
 sky130_fd_sc_hd__nor2_1 _1937_ (.A(_0319_),
    .B(_0337_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_0 _1938_ (.A1(_0313_),
    .A2(_0339_),
    .B1(\transfer_count[2][7] ),
    .Y(_0340_));
 sky130_fd_sc_hd__o31ai_1 _1939_ (.A1(\transfer_count[2][7] ),
    .A2(_0304_),
    .A3(_0338_),
    .B1(_0340_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand3_1 _1940_ (.A(\transfer_count[2][6] ),
    .B(\transfer_count[2][7] ),
    .C(_0331_),
    .Y(_0341_));
 sky130_fd_sc_hd__and2_0 _1941_ (.A(_0306_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__o21ai_0 _1942_ (.A1(_0313_),
    .A2(_0342_),
    .B1(\transfer_count[2][8] ),
    .Y(_0343_));
 sky130_fd_sc_hd__o31ai_1 _1943_ (.A1(\transfer_count[2][8] ),
    .A2(_0304_),
    .A3(_0341_),
    .B1(_0343_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand3_1 _1944_ (.A(\transfer_count[2][7] ),
    .B(\transfer_count[2][8] ),
    .C(_0337_),
    .Y(_0344_));
 sky130_fd_sc_hd__xor2_2 _1945_ (.A(\transfer_count[2][9] ),
    .B(_0344_),
    .X(_1375_));
 sky130_fd_sc_hd__and2_0 _1946_ (.A(_0306_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__o21ai_0 _1947_ (.A1(_0313_),
    .A2(_0345_),
    .B1(\transfer_count[2][9] ),
    .Y(_0346_));
 sky130_fd_sc_hd__o31ai_1 _1948_ (.A1(\transfer_count[2][9] ),
    .A2(_0304_),
    .A3(_0344_),
    .B1(_0346_),
    .Y(_0108_));
 sky130_fd_sc_hd__clkbuf_2 _1949_ (.A(\transfer_count[2][10] ),
    .X(_0347_));
 sky130_fd_sc_hd__and3_2 _1950_ (.A(\transfer_count[2][7] ),
    .B(\transfer_count[2][8] ),
    .C(\transfer_count[2][9] ),
    .X(_0348_));
 sky130_fd_sc_hd__nand4_4 _1951_ (.A(_0324_),
    .B(_0325_),
    .C(_0335_),
    .D(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__and3_1 _1952_ (.A(net140),
    .B(_0302_),
    .C(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__o21ai_0 _1953_ (.A1(_0313_),
    .A2(_0350_),
    .B1(_0347_),
    .Y(_0351_));
 sky130_fd_sc_hd__o31ai_1 _1954_ (.A1(_0347_),
    .A2(_0304_),
    .A3(_0349_),
    .B1(_0351_),
    .Y(_0078_));
 sky130_fd_sc_hd__nand3_1 _1955_ (.A(_0347_),
    .B(_0337_),
    .C(_0348_),
    .Y(_0352_));
 sky130_fd_sc_hd__xor2_1 _1956_ (.A(\transfer_count[2][11] ),
    .B(_0352_),
    .X(_1369_));
 sky130_fd_sc_hd__buf_2 _1957_ (.A(_0312_),
    .X(_0353_));
 sky130_fd_sc_hd__and2_0 _1958_ (.A(_0306_),
    .B(_0352_),
    .X(_0354_));
 sky130_fd_sc_hd__o21ai_0 _1959_ (.A1(_0353_),
    .A2(_0354_),
    .B1(\transfer_count[2][11] ),
    .Y(_0355_));
 sky130_fd_sc_hd__o31ai_1 _1960_ (.A1(\transfer_count[2][11] ),
    .A2(_0304_),
    .A3(_0352_),
    .B1(_0355_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(_0347_),
    .B(\transfer_count[2][11] ),
    .Y(_0356_));
 sky130_fd_sc_hd__nor2_1 _1962_ (.A(_0349_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_1 _1963_ (.A(_0316_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_1 _1964_ (.A(_0319_),
    .B(_0357_),
    .Y(_0359_));
 sky130_fd_sc_hd__o21ai_0 _1965_ (.A1(_0318_),
    .A2(_0359_),
    .B1(\transfer_count[2][12] ),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_0 _1966_ (.A1(\transfer_count[2][12] ),
    .A2(_0358_),
    .B1(_0360_),
    .Y(_0080_));
 sky130_fd_sc_hd__and2_0 _1967_ (.A(\transfer_count[2][11] ),
    .B(\transfer_count[2][12] ),
    .X(_0361_));
 sky130_fd_sc_hd__nand4_1 _1968_ (.A(_0347_),
    .B(_0337_),
    .C(_0348_),
    .D(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__xor2_1 _1969_ (.A(\transfer_count[2][13] ),
    .B(_0362_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_4 _1970_ (.A(_0303_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_0 _1971_ (.A(_0306_),
    .B(_0362_),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_0 _1972_ (.A1(_0353_),
    .A2(_0364_),
    .B1(\transfer_count[2][13] ),
    .Y(_0365_));
 sky130_fd_sc_hd__o31ai_1 _1973_ (.A1(\transfer_count[2][13] ),
    .A2(_0363_),
    .A3(_0362_),
    .B1(_0365_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand3_1 _1974_ (.A(\transfer_count[2][12] ),
    .B(\transfer_count[2][13] ),
    .C(_0357_),
    .Y(_0366_));
 sky130_fd_sc_hd__buf_2 _1975_ (.A(_0303_),
    .X(_0367_));
 sky130_fd_sc_hd__a31oi_1 _1976_ (.A1(\transfer_count[2][12] ),
    .A2(\transfer_count[2][13] ),
    .A3(_0357_),
    .B1(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21ai_0 _1977_ (.A1(_0353_),
    .A2(_0368_),
    .B1(\transfer_count[2][14] ),
    .Y(_0369_));
 sky130_fd_sc_hd__o31ai_1 _1978_ (.A1(\transfer_count[2][14] ),
    .A2(_0363_),
    .A3(_0366_),
    .B1(_0369_),
    .Y(_0082_));
 sky130_fd_sc_hd__clkbuf_2 _1979_ (.A(\transfer_count[2][15] ),
    .X(_0370_));
 sky130_fd_sc_hd__and3_1 _1980_ (.A(\transfer_count[2][12] ),
    .B(\transfer_count[2][13] ),
    .C(\transfer_count[2][14] ),
    .X(_0371_));
 sky130_fd_sc_hd__nand4_2 _1981_ (.A(_0347_),
    .B(\transfer_count[2][11] ),
    .C(_0348_),
    .D(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_4 _1982_ (.A(_0338_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__xnor2_1 _1983_ (.A(_0370_),
    .B(_0373_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _1984_ (.A(_0316_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__nor2_1 _1985_ (.A(_0367_),
    .B(_0373_),
    .Y(_0375_));
 sky130_fd_sc_hd__o21ai_0 _1986_ (.A1(_0318_),
    .A2(_0375_),
    .B1(_0370_),
    .Y(_0376_));
 sky130_fd_sc_hd__o21ai_0 _1987_ (.A1(_0370_),
    .A2(_0374_),
    .B1(_0376_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand3_1 _1988_ (.A(_0347_),
    .B(\transfer_count[2][11] ),
    .C(_0371_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _1989_ (.A(_0349_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__buf_2 _1990_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _1991_ (.A(_0370_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__a21oi_1 _1992_ (.A1(_0370_),
    .A2(_0379_),
    .B1(_0319_),
    .Y(_0381_));
 sky130_fd_sc_hd__o21ai_0 _1993_ (.A1(_0353_),
    .A2(_0381_),
    .B1(\transfer_count[2][16] ),
    .Y(_0382_));
 sky130_fd_sc_hd__o31ai_1 _1994_ (.A1(\transfer_count[2][16] ),
    .A2(_0363_),
    .A3(_0380_),
    .B1(_0382_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand3_1 _1995_ (.A(_0370_),
    .B(\transfer_count[2][16] ),
    .C(_0373_),
    .Y(_0383_));
 sky130_fd_sc_hd__a31oi_1 _1996_ (.A1(_0370_),
    .A2(\transfer_count[2][16] ),
    .A3(_0373_),
    .B1(_0367_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ai_0 _1997_ (.A1(_0353_),
    .A2(_0384_),
    .B1(\transfer_count[2][17] ),
    .Y(_0385_));
 sky130_fd_sc_hd__o31ai_1 _1998_ (.A1(\transfer_count[2][17] ),
    .A2(_0363_),
    .A3(_0383_),
    .B1(_0385_),
    .Y(_0085_));
 sky130_fd_sc_hd__and3_1 _1999_ (.A(_0370_),
    .B(\transfer_count[2][16] ),
    .C(\transfer_count[2][17] ),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_2 _2000_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _2001_ (.A(_0379_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _2002_ (.A1(_0379_),
    .A2(_0387_),
    .B1(_0319_),
    .Y(_0389_));
 sky130_fd_sc_hd__o21ai_0 _2003_ (.A1(_0353_),
    .A2(_0389_),
    .B1(\transfer_count[2][18] ),
    .Y(_0390_));
 sky130_fd_sc_hd__o31ai_1 _2004_ (.A1(\transfer_count[2][18] ),
    .A2(_0363_),
    .A3(_0388_),
    .B1(_0390_),
    .Y(_0086_));
 sky130_fd_sc_hd__nand3_1 _2005_ (.A(\transfer_count[2][18] ),
    .B(_0373_),
    .C(_0387_),
    .Y(_0391_));
 sky130_fd_sc_hd__xor2_1 _2006_ (.A(\transfer_count[2][19] ),
    .B(_0391_),
    .X(_1345_));
 sky130_fd_sc_hd__a31oi_1 _2007_ (.A1(\transfer_count[2][18] ),
    .A2(_0373_),
    .A3(_0387_),
    .B1(_0367_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_0 _2008_ (.A1(_0353_),
    .A2(_0392_),
    .B1(\transfer_count[2][19] ),
    .Y(_0393_));
 sky130_fd_sc_hd__o31ai_1 _2009_ (.A1(\transfer_count[2][19] ),
    .A2(_0363_),
    .A3(_0391_),
    .B1(_0393_),
    .Y(_0087_));
 sky130_fd_sc_hd__nand3_1 _2010_ (.A(_0370_),
    .B(\transfer_count[2][16] ),
    .C(\transfer_count[2][17] ),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_1 _2011_ (.A(\transfer_count[2][18] ),
    .B(\transfer_count[2][19] ),
    .Y(_0395_));
 sky130_fd_sc_hd__nor4_1 _2012_ (.A(_0349_),
    .B(_0377_),
    .C(_0394_),
    .D(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nand2_1 _2013_ (.A(_0316_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__nor2_1 _2014_ (.A(_0367_),
    .B(_0396_),
    .Y(_0398_));
 sky130_fd_sc_hd__o21ai_0 _2015_ (.A1(_0318_),
    .A2(_0398_),
    .B1(\transfer_count[2][20] ),
    .Y(_0399_));
 sky130_fd_sc_hd__o21ai_0 _2016_ (.A1(\transfer_count[2][20] ),
    .A2(_0397_),
    .B1(_0399_),
    .Y(_0089_));
 sky130_fd_sc_hd__and3_1 _2017_ (.A(\transfer_count[2][18] ),
    .B(\transfer_count[2][19] ),
    .C(\transfer_count[2][20] ),
    .X(_0400_));
 sky130_fd_sc_hd__nand3_1 _2018_ (.A(_0373_),
    .B(_0387_),
    .C(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xor2_1 _2019_ (.A(\transfer_count[2][21] ),
    .B(_0401_),
    .X(_1339_));
 sky130_fd_sc_hd__a31oi_1 _2020_ (.A1(_0373_),
    .A2(_0387_),
    .A3(_0400_),
    .B1(_0367_),
    .Y(_0402_));
 sky130_fd_sc_hd__o21ai_0 _2021_ (.A1(_0353_),
    .A2(_0402_),
    .B1(\transfer_count[2][21] ),
    .Y(_0403_));
 sky130_fd_sc_hd__o31ai_1 _2022_ (.A1(\transfer_count[2][21] ),
    .A2(_0363_),
    .A3(_0401_),
    .B1(_0403_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_1 _2023_ (.A(\transfer_count[2][22] ),
    .Y(_0404_));
 sky130_fd_sc_hd__nand4_1 _2024_ (.A(\transfer_count[2][21] ),
    .B(_0378_),
    .C(_0387_),
    .D(_0400_),
    .Y(_0405_));
 sky130_fd_sc_hd__a21oi_1 _2025_ (.A1(_0316_),
    .A2(_0405_),
    .B1(_0312_),
    .Y(_0406_));
 sky130_fd_sc_hd__or3_1 _2026_ (.A(\transfer_count[2][22] ),
    .B(_0303_),
    .C(_0405_),
    .X(_0407_));
 sky130_fd_sc_hd__o21ai_0 _2027_ (.A1(_0404_),
    .A2(_0406_),
    .B1(_0407_),
    .Y(_0091_));
 sky130_fd_sc_hd__clkbuf_2 _2028_ (.A(\transfer_count[2][23] ),
    .X(_0408_));
 sky130_fd_sc_hd__and4_1 _2029_ (.A(\transfer_count[2][21] ),
    .B(\transfer_count[2][22] ),
    .C(_0387_),
    .D(_0400_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_2 _2030_ (.A(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__nor3b_1 _2031_ (.A(_0338_),
    .B(_0372_),
    .C_N(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__buf_2 _2032_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__xnor2_1 _2033_ (.A(_0408_),
    .B(_0412_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _2034_ (.A(_0316_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__nor2_1 _2035_ (.A(_0367_),
    .B(_0412_),
    .Y(_0414_));
 sky130_fd_sc_hd__o21ai_0 _2036_ (.A1(_0318_),
    .A2(_0414_),
    .B1(_0408_),
    .Y(_0415_));
 sky130_fd_sc_hd__o21ai_0 _2037_ (.A1(_0408_),
    .A2(_0413_),
    .B1(_0415_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand3_1 _2038_ (.A(_0408_),
    .B(_0379_),
    .C(_0410_),
    .Y(_0416_));
 sky130_fd_sc_hd__a31oi_1 _2039_ (.A1(_0408_),
    .A2(_0379_),
    .A3(_0410_),
    .B1(_0367_),
    .Y(_0417_));
 sky130_fd_sc_hd__o21ai_0 _2040_ (.A1(_0353_),
    .A2(_0417_),
    .B1(\transfer_count[2][24] ),
    .Y(_0418_));
 sky130_fd_sc_hd__o31ai_1 _2041_ (.A1(\transfer_count[2][24] ),
    .A2(_0363_),
    .A3(_0416_),
    .B1(_0418_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand3_1 _2042_ (.A(_0408_),
    .B(\transfer_count[2][24] ),
    .C(_0412_),
    .Y(_0419_));
 sky130_fd_sc_hd__xor2_1 _2043_ (.A(\transfer_count[2][25] ),
    .B(_0419_),
    .X(_1327_));
 sky130_fd_sc_hd__a31oi_1 _2044_ (.A1(_0408_),
    .A2(\transfer_count[2][24] ),
    .A3(_0412_),
    .B1(_0367_),
    .Y(_0420_));
 sky130_fd_sc_hd__o21ai_0 _2045_ (.A1(_0353_),
    .A2(_0420_),
    .B1(\transfer_count[2][25] ),
    .Y(_0421_));
 sky130_fd_sc_hd__o31ai_1 _2046_ (.A1(\transfer_count[2][25] ),
    .A2(_0363_),
    .A3(_0419_),
    .B1(_0421_),
    .Y(_0094_));
 sky130_fd_sc_hd__and3_1 _2047_ (.A(_0408_),
    .B(\transfer_count[2][24] ),
    .C(\transfer_count[2][25] ),
    .X(_0422_));
 sky130_fd_sc_hd__nand3_1 _2048_ (.A(_0379_),
    .B(_0410_),
    .C(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a31oi_1 _2049_ (.A1(_0379_),
    .A2(_0410_),
    .A3(_0422_),
    .B1(_0367_),
    .Y(_0424_));
 sky130_fd_sc_hd__o21ai_0 _2050_ (.A1(_0318_),
    .A2(_0424_),
    .B1(\transfer_count[2][26] ),
    .Y(_0425_));
 sky130_fd_sc_hd__o31ai_1 _2051_ (.A1(\transfer_count[2][26] ),
    .A2(_0363_),
    .A3(_0423_),
    .B1(_0425_),
    .Y(_0095_));
 sky130_fd_sc_hd__and3_1 _2052_ (.A(\transfer_count[2][26] ),
    .B(_0411_),
    .C(_0422_),
    .X(_0426_));
 sky130_fd_sc_hd__xnor2_1 _2053_ (.A(\transfer_count[2][27] ),
    .B(_0426_),
    .Y(_1321_));
 sky130_fd_sc_hd__nand2_1 _2054_ (.A(_0316_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__a31oi_1 _2055_ (.A1(\transfer_count[2][26] ),
    .A2(_0412_),
    .A3(_0422_),
    .B1(_0303_),
    .Y(_0428_));
 sky130_fd_sc_hd__o21ai_0 _2056_ (.A1(_0312_),
    .A2(_0428_),
    .B1(\transfer_count[2][27] ),
    .Y(_0429_));
 sky130_fd_sc_hd__o21ai_0 _2057_ (.A1(\transfer_count[2][27] ),
    .A2(_0427_),
    .B1(_0429_),
    .Y(_0096_));
 sky130_fd_sc_hd__and3_1 _2058_ (.A(\transfer_count[2][26] ),
    .B(\transfer_count[2][27] ),
    .C(_0422_),
    .X(_0430_));
 sky130_fd_sc_hd__nand3_1 _2059_ (.A(_0379_),
    .B(_0410_),
    .C(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a31oi_1 _2060_ (.A1(_0379_),
    .A2(_0410_),
    .A3(_0430_),
    .B1(_0303_),
    .Y(_0432_));
 sky130_fd_sc_hd__o21ai_0 _2061_ (.A1(_0318_),
    .A2(_0432_),
    .B1(\transfer_count[2][28] ),
    .Y(_0433_));
 sky130_fd_sc_hd__o31ai_1 _2062_ (.A1(\transfer_count[2][28] ),
    .A2(_0319_),
    .A3(_0431_),
    .B1(_0433_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand3_1 _2063_ (.A(\transfer_count[2][28] ),
    .B(_0412_),
    .C(_0430_),
    .Y(_0434_));
 sky130_fd_sc_hd__xor2_1 _2064_ (.A(\transfer_count[2][29] ),
    .B(_0434_),
    .X(_1315_));
 sky130_fd_sc_hd__a31oi_1 _2065_ (.A1(\transfer_count[2][28] ),
    .A2(_0412_),
    .A3(_0430_),
    .B1(_0303_),
    .Y(_0435_));
 sky130_fd_sc_hd__o21ai_0 _2066_ (.A1(_0318_),
    .A2(_0435_),
    .B1(\transfer_count[2][29] ),
    .Y(_0436_));
 sky130_fd_sc_hd__o31ai_1 _2067_ (.A1(\transfer_count[2][29] ),
    .A2(_0319_),
    .A3(_0434_),
    .B1(_0436_),
    .Y(_0098_));
 sky130_fd_sc_hd__and3_1 _2068_ (.A(\transfer_count[2][28] ),
    .B(\transfer_count[2][29] ),
    .C(_0430_),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _2069_ (.A(_0378_),
    .B(_0410_),
    .C(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__nand2b_1 _2070_ (.A_N(_0438_),
    .B(_0306_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor2b_1 _2071_ (.A(_0312_),
    .B_N(\transfer_count[2][30] ),
    .Y(_0440_));
 sky130_fd_sc_hd__a21oi_1 _2072_ (.A1(_0316_),
    .A2(_0438_),
    .B1(\transfer_count[2][30] ),
    .Y(_0441_));
 sky130_fd_sc_hd__a21oi_1 _2073_ (.A1(_0439_),
    .A2(_0440_),
    .B1(_0441_),
    .Y(_0100_));
 sky130_fd_sc_hd__nand3_1 _2074_ (.A(\transfer_count[2][30] ),
    .B(_0412_),
    .C(_0437_),
    .Y(_0442_));
 sky130_fd_sc_hd__a31oi_1 _2075_ (.A1(\transfer_count[2][30] ),
    .A2(_0412_),
    .A3(_0437_),
    .B1(_0303_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21ai_0 _2076_ (.A1(_0318_),
    .A2(_0443_),
    .B1(\transfer_count[2][31] ),
    .Y(_0444_));
 sky130_fd_sc_hd__o31ai_1 _2077_ (.A1(\transfer_count[2][31] ),
    .A2(_0319_),
    .A3(_0442_),
    .B1(_0444_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_1 _2078_ (.A(\transfer_count[1][0] ),
    .Y(_1409_));
 sky130_fd_sc_hd__buf_2 _2079_ (.A(\channel_state[1][2] ),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_2 _2080_ (.A(net139),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21boi_4 _2081_ (.A1(_0446_),
    .A2(_0882_),
    .B1_N(_0827_),
    .Y(_0447_));
 sky130_fd_sc_hd__clkbuf_4 _2082_ (.A(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__nor3_4 _2083_ (.A(_0825_),
    .B(_0826_),
    .C(_0446_),
    .Y(_0449_));
 sky130_fd_sc_hd__clkbuf_4 _2084_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _2085_ (.A(\transfer_count[1][0] ),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__a21oi_1 _2086_ (.A1(\transfer_count[1][0] ),
    .A2(_0448_),
    .B1(_0451_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _2087_ (.A(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__buf_2 _2088_ (.A(_0828_),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _2089_ (.A(_0446_),
    .B(_0882_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_4 _2090_ (.A(_0827_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__clkbuf_4 _2091_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _2092_ (.A(\transfer_count[1][1] ),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_0 _2093_ (.A1(_1414_),
    .A2(_0452_),
    .B1(_0456_),
    .Y(_0056_));
 sky130_fd_sc_hd__nand2_1 _2094_ (.A(_1412_),
    .B(_0450_),
    .Y(_0457_));
 sky130_fd_sc_hd__o21ai_0 _2095_ (.A1(_1412_),
    .A2(_0828_),
    .B1(_0447_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _2096_ (.A(\transfer_count[1][2] ),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__o21ai_0 _2097_ (.A1(\transfer_count[1][2] ),
    .A2(_0457_),
    .B1(_0459_),
    .Y(_0067_));
 sky130_fd_sc_hd__nand3_1 _2098_ (.A(\transfer_count[1][0] ),
    .B(\transfer_count[1][1] ),
    .C(\transfer_count[1][2] ),
    .Y(_0460_));
 sky130_fd_sc_hd__and2_0 _2099_ (.A(_0449_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__o21ai_0 _2100_ (.A1(_0454_),
    .A2(_0461_),
    .B1(\transfer_count[1][3] ),
    .Y(_0462_));
 sky130_fd_sc_hd__o31ai_1 _2101_ (.A1(\transfer_count[1][3] ),
    .A2(_0829_),
    .A3(_0460_),
    .B1(_0462_),
    .Y(_0070_));
 sky130_fd_sc_hd__nand3_2 _2102_ (.A(_1412_),
    .B(\transfer_count[1][2] ),
    .C(\transfer_count[1][3] ),
    .Y(_0463_));
 sky130_fd_sc_hd__xor2_1 _2103_ (.A(\transfer_count[1][4] ),
    .B(_0463_),
    .X(_1432_));
 sky130_fd_sc_hd__nand2_1 _2104_ (.A(\transfer_count[1][4] ),
    .B(_0455_),
    .Y(_0464_));
 sky130_fd_sc_hd__o21ai_0 _2105_ (.A1(_0452_),
    .A2(_1432_),
    .B1(_0464_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(\transfer_count[1][3] ),
    .B(\transfer_count[1][4] ),
    .Y(_0465_));
 sky130_fd_sc_hd__nor2_1 _2107_ (.A(_0460_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__xnor2_1 _2108_ (.A(\transfer_count[1][5] ),
    .B(_0466_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _2109_ (.A(\transfer_count[1][5] ),
    .B(_0455_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_0 _2110_ (.A1(_0452_),
    .A2(_1429_),
    .B1(_0467_),
    .Y(_0072_));
 sky130_fd_sc_hd__nor2_1 _2111_ (.A(_0798_),
    .B(_0463_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _2112_ (.A(_0450_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21ai_0 _2113_ (.A1(_0828_),
    .A2(_0468_),
    .B1(_0447_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _2114_ (.A(_0800_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__o21ai_0 _2115_ (.A1(_0800_),
    .A2(_0469_),
    .B1(_0471_),
    .Y(_0073_));
 sky130_fd_sc_hd__nor3_1 _2116_ (.A(_0797_),
    .B(_0798_),
    .C(_0799_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _2117_ (.A(_0800_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a21oi_1 _2118_ (.A1(_0800_),
    .A2(_0472_),
    .B1(_0829_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_0 _2119_ (.A1(_0454_),
    .A2(_0474_),
    .B1(\transfer_count[1][7] ),
    .Y(_0475_));
 sky130_fd_sc_hd__o31ai_1 _2120_ (.A1(\transfer_count[1][7] ),
    .A2(_0829_),
    .A3(_0473_),
    .B1(_0475_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand3_1 _2121_ (.A(\transfer_count[1][7] ),
    .B(_0800_),
    .C(_0468_),
    .Y(_0476_));
 sky130_fd_sc_hd__nor3_4 _2122_ (.A(_0798_),
    .B(_0801_),
    .C(_0463_),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_0 _2123_ (.A1(_0829_),
    .A2(_0477_),
    .B1(_0447_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _2124_ (.A(\transfer_count[1][8] ),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o31ai_1 _2125_ (.A1(\transfer_count[1][8] ),
    .A2(_0829_),
    .A3(_0476_),
    .B1(_0479_),
    .Y(_0075_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(\transfer_count[1][9] ),
    .B(_0455_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_0 _2127_ (.A1(_1051_),
    .A2(_0452_),
    .B1(_0480_),
    .Y(_0076_));
 sky130_fd_sc_hd__and3_1 _2128_ (.A(\transfer_count[1][9] ),
    .B(\transfer_count[1][8] ),
    .C(_0477_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_1 _2129_ (.A(\transfer_count[1][10] ),
    .B(_0481_),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _2130_ (.A(\transfer_count[1][10] ),
    .B(_0455_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ai_0 _2131_ (.A1(_0452_),
    .A2(_1048_),
    .B1(_0482_),
    .Y(_0046_));
 sky130_fd_sc_hd__nand2_1 _2132_ (.A(_0803_),
    .B(_0804_),
    .Y(_0483_));
 sky130_fd_sc_hd__xor2_1 _2133_ (.A(\transfer_count[1][11] ),
    .B(_0483_),
    .X(_1045_));
 sky130_fd_sc_hd__nand2_1 _2134_ (.A(\transfer_count[1][11] ),
    .B(_0455_),
    .Y(_0484_));
 sky130_fd_sc_hd__o21ai_0 _2135_ (.A1(_0452_),
    .A2(_1045_),
    .B1(_0484_),
    .Y(_0047_));
 sky130_fd_sc_hd__and3_1 _2136_ (.A(\transfer_count[1][11] ),
    .B(_0804_),
    .C(_0477_),
    .X(_0485_));
 sky130_fd_sc_hd__xnor2_1 _2137_ (.A(\transfer_count[1][12] ),
    .B(_0485_),
    .Y(_1042_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(\transfer_count[1][12] ),
    .B(_0455_),
    .Y(_0486_));
 sky130_fd_sc_hd__o21ai_0 _2139_ (.A1(_0452_),
    .A2(_1042_),
    .B1(_0486_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _2140_ (.A(_0805_),
    .B(_0450_),
    .Y(_0487_));
 sky130_fd_sc_hd__o21ai_0 _2141_ (.A1(_0805_),
    .A2(_0828_),
    .B1(_0447_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _2142_ (.A(\transfer_count[1][13] ),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_0 _2143_ (.A1(\transfer_count[1][13] ),
    .A2(_0487_),
    .B1(_0489_),
    .Y(_0049_));
 sky130_fd_sc_hd__or2_0 _2144_ (.A(_0809_),
    .B(_0810_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_1 _2145_ (.A(_0490_),
    .B(_0476_),
    .Y(_0491_));
 sky130_fd_sc_hd__xnor2_1 _2146_ (.A(\transfer_count[1][14] ),
    .B(_0491_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand2_1 _2147_ (.A(\transfer_count[1][14] ),
    .B(_0455_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21ai_0 _2148_ (.A1(_0452_),
    .A2(_1036_),
    .B1(_0492_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_1 _2149_ (.A(_0490_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand3_1 _2150_ (.A(\transfer_count[1][14] ),
    .B(_0803_),
    .C(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__xor2_1 _2151_ (.A(\transfer_count[1][15] ),
    .B(_0494_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _2152_ (.A(\transfer_count[1][15] ),
    .B(_0455_),
    .Y(_0495_));
 sky130_fd_sc_hd__o21ai_0 _2153_ (.A1(_0452_),
    .A2(_1033_),
    .B1(_0495_),
    .Y(_0051_));
 sky130_fd_sc_hd__nor3b_1 _2154_ (.A(_0490_),
    .B(_0811_),
    .C_N(_0477_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _2155_ (.A(_0450_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__o21ai_0 _2156_ (.A1(_0828_),
    .A2(_0496_),
    .B1(_0447_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_1 _2157_ (.A(\transfer_count[1][16] ),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21ai_0 _2158_ (.A1(\transfer_count[1][16] ),
    .A2(_0497_),
    .B1(_0499_),
    .Y(_0052_));
 sky130_fd_sc_hd__a21oi_1 _2159_ (.A1(_0803_),
    .A2(_0812_),
    .B1(_0829_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_0 _2160_ (.A1(_0454_),
    .A2(_0500_),
    .B1(_0813_),
    .Y(_0501_));
 sky130_fd_sc_hd__o31ai_1 _2161_ (.A1(_0813_),
    .A2(_0823_),
    .A3(_0829_),
    .B1(_0501_),
    .Y(_0053_));
 sky130_fd_sc_hd__and2_0 _2162_ (.A(_0812_),
    .B(_0477_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_2 _2163_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_1 _2164_ (.A(_0813_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _2165_ (.A(_0450_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a31oi_1 _2166_ (.A1(_0813_),
    .A2(_0449_),
    .A3(_0503_),
    .B1(\transfer_count[1][18] ),
    .Y(_0506_));
 sky130_fd_sc_hd__a31oi_1 _2167_ (.A1(\transfer_count[1][18] ),
    .A2(_0448_),
    .A3(_0505_),
    .B1(_0506_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _2168_ (.A(\transfer_count[1][18] ),
    .B(_0813_),
    .Y(_0507_));
 sky130_fd_sc_hd__buf_2 _2169_ (.A(_0449_),
    .X(_0508_));
 sky130_fd_sc_hd__o21ai_0 _2170_ (.A1(_0507_),
    .A2(_0823_),
    .B1(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nor2_1 _2171_ (.A(_0507_),
    .B(_0823_),
    .Y(_0510_));
 sky130_fd_sc_hd__a21oi_1 _2172_ (.A1(_0510_),
    .A2(_0508_),
    .B1(\transfer_count[1][19] ),
    .Y(_0511_));
 sky130_fd_sc_hd__a31oi_1 _2173_ (.A1(\transfer_count[1][19] ),
    .A2(_0448_),
    .A3(_0509_),
    .B1(_0511_),
    .Y(_0055_));
 sky130_fd_sc_hd__and3_1 _2174_ (.A(\transfer_count[1][19] ),
    .B(\transfer_count[1][18] ),
    .C(_0813_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _2175_ (.A(_0512_),
    .B(_0503_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _2176_ (.A(_0450_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__a31oi_1 _2177_ (.A1(_0512_),
    .A2(_0449_),
    .A3(_0503_),
    .B1(\transfer_count[1][20] ),
    .Y(_0515_));
 sky130_fd_sc_hd__a31oi_1 _2178_ (.A1(\transfer_count[1][20] ),
    .A2(_0448_),
    .A3(_0514_),
    .B1(_0515_),
    .Y(_0057_));
 sky130_fd_sc_hd__o21ai_0 _2179_ (.A1(_0814_),
    .A2(_0823_),
    .B1(_0508_),
    .Y(_0516_));
 sky130_fd_sc_hd__a21oi_1 _2180_ (.A1(_0824_),
    .A2(_0508_),
    .B1(\transfer_count[1][21] ),
    .Y(_0517_));
 sky130_fd_sc_hd__a31oi_1 _2181_ (.A1(\transfer_count[1][21] ),
    .A2(_0448_),
    .A3(_0516_),
    .B1(_0517_),
    .Y(_0058_));
 sky130_fd_sc_hd__and3_1 _2182_ (.A(\transfer_count[1][21] ),
    .B(\transfer_count[1][20] ),
    .C(_0512_),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _2183_ (.A(_0518_),
    .B(_0503_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _2184_ (.A(_0450_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a31oi_1 _2185_ (.A1(_0518_),
    .A2(_0449_),
    .A3(_0503_),
    .B1(\transfer_count[1][22] ),
    .Y(_0521_));
 sky130_fd_sc_hd__a31oi_1 _2186_ (.A1(\transfer_count[1][22] ),
    .A2(_0448_),
    .A3(_0520_),
    .B1(_0521_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand2_1 _2187_ (.A(_0803_),
    .B(_0818_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _2188_ (.A(_0522_),
    .B(_0508_),
    .Y(_0523_));
 sky130_fd_sc_hd__a31oi_1 _2189_ (.A1(_0803_),
    .A2(_0818_),
    .A3(_0449_),
    .B1(\transfer_count[1][23] ),
    .Y(_0524_));
 sky130_fd_sc_hd__a31oi_1 _2190_ (.A1(\transfer_count[1][23] ),
    .A2(_0448_),
    .A3(_0523_),
    .B1(_0524_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand3_1 _2191_ (.A(\transfer_count[1][23] ),
    .B(_0818_),
    .C(_0477_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _2192_ (.A(_0450_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__a41oi_1 _2193_ (.A1(\transfer_count[1][23] ),
    .A2(_0818_),
    .A3(_0449_),
    .A4(_0477_),
    .B1(\transfer_count[1][24] ),
    .Y(_0527_));
 sky130_fd_sc_hd__a31oi_1 _2194_ (.A1(\transfer_count[1][24] ),
    .A2(_0448_),
    .A3(_0526_),
    .B1(_0527_),
    .Y(_0061_));
 sky130_fd_sc_hd__a21oi_1 _2195_ (.A1(_0822_),
    .A2(_0449_),
    .B1(_0454_),
    .Y(_0528_));
 sky130_fd_sc_hd__or3_1 _2196_ (.A(\transfer_count[1][25] ),
    .B(_0822_),
    .C(_0828_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_0 _2197_ (.A1(_0821_),
    .A2(_0528_),
    .B1(_0529_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand4_2 _2198_ (.A(_0812_),
    .B(_0816_),
    .C(_0819_),
    .D(_0477_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _2199_ (.A(_0450_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nor2_1 _2200_ (.A(_0829_),
    .B(_0530_),
    .Y(_0532_));
 sky130_fd_sc_hd__nor2_1 _2201_ (.A(\transfer_count[1][26] ),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a31oi_1 _2202_ (.A1(\transfer_count[1][26] ),
    .A2(_0448_),
    .A3(_0531_),
    .B1(_0533_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_1 _2203_ (.A(\transfer_count[1][27] ),
    .Y(_0534_));
 sky130_fd_sc_hd__nand4_1 _2204_ (.A(\transfer_count[1][26] ),
    .B(_0803_),
    .C(_0818_),
    .D(_0819_),
    .Y(_0535_));
 sky130_fd_sc_hd__a21oi_1 _2205_ (.A1(_0449_),
    .A2(_0535_),
    .B1(_0454_),
    .Y(_0536_));
 sky130_fd_sc_hd__or3_1 _2206_ (.A(\transfer_count[1][27] ),
    .B(_0828_),
    .C(_0535_),
    .X(_0537_));
 sky130_fd_sc_hd__o21ai_0 _2207_ (.A1(_0534_),
    .A2(_0536_),
    .B1(_0537_),
    .Y(_0064_));
 sky130_fd_sc_hd__nand2_1 _2208_ (.A(\transfer_count[1][27] ),
    .B(\transfer_count[1][26] ),
    .Y(_0538_));
 sky130_fd_sc_hd__o21ai_0 _2209_ (.A1(_0538_),
    .A2(_0530_),
    .B1(_0508_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_1 _2210_ (.A(_0538_),
    .B(_0530_),
    .Y(_0540_));
 sky130_fd_sc_hd__a21oi_1 _2211_ (.A1(_0508_),
    .A2(_0540_),
    .B1(\transfer_count[1][28] ),
    .Y(_0541_));
 sky130_fd_sc_hd__a31oi_1 _2212_ (.A1(\transfer_count[1][28] ),
    .A2(_0448_),
    .A3(_0539_),
    .B1(_0541_),
    .Y(_0065_));
 sky130_fd_sc_hd__nand2_1 _2213_ (.A(_0820_),
    .B(_0508_),
    .Y(_0542_));
 sky130_fd_sc_hd__o21ba_1 _2214_ (.A1(_0820_),
    .A2(_0828_),
    .B1_N(\transfer_count[1][29] ),
    .X(_0543_));
 sky130_fd_sc_hd__a31oi_1 _2215_ (.A1(\transfer_count[1][29] ),
    .A2(_0447_),
    .A3(_0542_),
    .B1(_0543_),
    .Y(_0066_));
 sky130_fd_sc_hd__and3_1 _2216_ (.A(\transfer_count[1][29] ),
    .B(_0807_),
    .C(_0819_),
    .X(_0544_));
 sky130_fd_sc_hd__nand4_2 _2217_ (.A(_0812_),
    .B(_0816_),
    .C(_0477_),
    .D(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _2218_ (.A(_0508_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nor2_1 _2219_ (.A(_0829_),
    .B(_0545_),
    .Y(_0547_));
 sky130_fd_sc_hd__nor2_1 _2220_ (.A(\transfer_count[1][30] ),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a31oi_1 _2221_ (.A1(\transfer_count[1][30] ),
    .A2(_0447_),
    .A3(_0546_),
    .B1(_0548_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _2222_ (.A(\transfer_count[1][30] ),
    .B(\transfer_count[1][29] ),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_0 _2223_ (.A1(_0820_),
    .A2(_0549_),
    .B1(_0508_),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_1 _2224_ (.A(\transfer_count[1][31] ),
    .Y(_0551_));
 sky130_fd_sc_hd__o31a_1 _2225_ (.A1(_0820_),
    .A2(_0828_),
    .A3(_0549_),
    .B1(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a31oi_1 _2226_ (.A1(\transfer_count[1][31] ),
    .A2(_0447_),
    .A3(_0550_),
    .B1(_0552_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_1 _2227_ (.A(\transfer_count[0][0] ),
    .Y(_1205_));
 sky130_fd_sc_hd__buf_2 _2228_ (.A(\channel_state[0][2] ),
    .X(_0553_));
 sky130_fd_sc_hd__nor2_1 _2229_ (.A(_0980_),
    .B(_0981_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand3_2 _2230_ (.A(net138),
    .B(_0553_),
    .C(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__buf_2 _2231_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__nor2_2 _2232_ (.A(_0148_),
    .B(_0202_),
    .Y(_0557_));
 sky130_fd_sc_hd__clkbuf_4 _2233_ (.A(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _2234_ (.A(\transfer_count[0][0] ),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__o21ai_0 _2235_ (.A1(\transfer_count[0][0] ),
    .A2(_0556_),
    .B1(_0559_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_1 _2236_ (.A(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__clkbuf_4 _2237_ (.A(_0555_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(\transfer_count[0][1] ),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__o22ai_1 _2239_ (.A1(_1210_),
    .A2(_0556_),
    .B1(_0202_),
    .B2(_0561_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _2240_ (.A(_1208_),
    .B(_0150_),
    .Y(_0562_));
 sky130_fd_sc_hd__clkbuf_4 _2241_ (.A(_0557_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_4 _2242_ (.A(_0555_),
    .X(_0564_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_1208_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_0 _2244_ (.A1(_0563_),
    .A2(_0565_),
    .B1(\transfer_count[0][2] ),
    .Y(_0566_));
 sky130_fd_sc_hd__o21ai_0 _2245_ (.A1(\transfer_count[0][2] ),
    .A2(_0562_),
    .B1(_0566_),
    .Y(_0035_));
 sky130_fd_sc_hd__nand2_1 _2246_ (.A(_0987_),
    .B(_0150_),
    .Y(_0567_));
 sky130_fd_sc_hd__nor2_1 _2247_ (.A(_0987_),
    .B(_0564_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_0 _2248_ (.A1(_0557_),
    .A2(_0568_),
    .B1(\transfer_count[0][3] ),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_0 _2249_ (.A1(\transfer_count[0][3] ),
    .A2(_0567_),
    .B1(_0569_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand3_1 _2250_ (.A(\transfer_count[0][2] ),
    .B(\transfer_count[0][3] ),
    .C(_1208_),
    .Y(_0570_));
 sky130_fd_sc_hd__xor2_1 _2251_ (.A(\transfer_count[0][4] ),
    .B(_0570_),
    .X(_1228_));
 sky130_fd_sc_hd__nand2_1 _2252_ (.A(\transfer_count[0][4] ),
    .B(_0560_),
    .Y(_0571_));
 sky130_fd_sc_hd__o22ai_1 _2253_ (.A1(_0556_),
    .A2(_1228_),
    .B1(_0571_),
    .B2(_0202_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand2_1 _2254_ (.A(\transfer_count[0][5] ),
    .B(_0558_),
    .Y(_0572_));
 sky130_fd_sc_hd__o21ai_0 _2255_ (.A1(_1225_),
    .A2(_0556_),
    .B1(_0572_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand3_2 _2256_ (.A(\transfer_count[0][2] ),
    .B(_1208_),
    .C(_0992_),
    .Y(_0573_));
 sky130_fd_sc_hd__and2_0 _2257_ (.A(_0149_),
    .B(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__o21ai_0 _2258_ (.A1(_0558_),
    .A2(_0574_),
    .B1(\transfer_count[0][6] ),
    .Y(_0575_));
 sky130_fd_sc_hd__o31ai_1 _2259_ (.A1(\transfer_count[0][6] ),
    .A2(_0560_),
    .A3(_0573_),
    .B1(_0575_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _2260_ (.A(_0997_),
    .B(_0150_),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_1 _2261_ (.A(_0997_),
    .B(_0564_),
    .Y(_0577_));
 sky130_fd_sc_hd__o21ai_0 _2262_ (.A1(_0557_),
    .A2(_0577_),
    .B1(_0991_),
    .Y(_0578_));
 sky130_fd_sc_hd__o21ai_0 _2263_ (.A1(_0991_),
    .A2(_0576_),
    .B1(_0578_),
    .Y(_0042_));
 sky130_fd_sc_hd__and2_0 _2264_ (.A(\transfer_count[0][6] ),
    .B(_0991_),
    .X(_0579_));
 sky130_fd_sc_hd__nand4_4 _2265_ (.A(\transfer_count[0][2] ),
    .B(_1208_),
    .C(_0992_),
    .D(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2b_1 _2266_ (.A(_0573_),
    .B_N(_0579_),
    .Y(_0581_));
 sky130_fd_sc_hd__nor2_1 _2267_ (.A(_0564_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__o21ai_0 _2268_ (.A1(_0558_),
    .A2(_0582_),
    .B1(_0989_),
    .Y(_0583_));
 sky130_fd_sc_hd__o31ai_1 _2269_ (.A1(_0989_),
    .A2(_0560_),
    .A3(_0580_),
    .B1(_0583_),
    .Y(_0043_));
 sky130_fd_sc_hd__clkbuf_4 _2270_ (.A(_0555_),
    .X(_0584_));
 sky130_fd_sc_hd__a31oi_1 _2271_ (.A1(_0991_),
    .A2(_0989_),
    .A3(_0997_),
    .B1(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o21ai_0 _2272_ (.A1(_0558_),
    .A2(_0585_),
    .B1(\transfer_count[0][9] ),
    .Y(_0586_));
 sky130_fd_sc_hd__o31ai_1 _2273_ (.A1(\transfer_count[0][9] ),
    .A2(_0998_),
    .A3(_0556_),
    .B1(_0586_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand3_1 _2274_ (.A(\transfer_count[0][9] ),
    .B(_0989_),
    .C(_0581_),
    .Y(_0587_));
 sky130_fd_sc_hd__xor2_1 _2275_ (.A(\transfer_count[0][10] ),
    .B(_0587_),
    .X(_1246_));
 sky130_fd_sc_hd__nand2_1 _2276_ (.A(\transfer_count[0][10] ),
    .B(_0558_),
    .Y(_0588_));
 sky130_fd_sc_hd__o21ai_0 _2277_ (.A1(_0556_),
    .A2(_1246_),
    .B1(_0588_),
    .Y(_0014_));
 sky130_fd_sc_hd__and3_1 _2278_ (.A(_0991_),
    .B(_1006_),
    .C(_0997_),
    .X(_0589_));
 sky130_fd_sc_hd__nand2_1 _2279_ (.A(_0589_),
    .B(_0150_),
    .Y(_0590_));
 sky130_fd_sc_hd__or2_0 _2280_ (.A(_0149_),
    .B(_0202_),
    .X(_0591_));
 sky130_fd_sc_hd__buf_2 _2281_ (.A(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__o21ai_0 _2282_ (.A1(_0994_),
    .A2(_0564_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _2283_ (.A(\transfer_count[0][11] ),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__o21ai_0 _2284_ (.A1(\transfer_count[0][11] ),
    .A2(_0590_),
    .B1(_0594_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand3_1 _2285_ (.A(\transfer_count[0][11] ),
    .B(_1006_),
    .C(_0581_),
    .Y(_0595_));
 sky130_fd_sc_hd__xor2_1 _2286_ (.A(\transfer_count[0][12] ),
    .B(_0595_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _2287_ (.A(\transfer_count[0][12] ),
    .B(_0558_),
    .Y(_0596_));
 sky130_fd_sc_hd__o21ai_0 _2288_ (.A1(_0556_),
    .A2(_1240_),
    .B1(_0596_),
    .Y(_0016_));
 sky130_fd_sc_hd__a31oi_1 _2289_ (.A1(\transfer_count[0][12] ),
    .A2(\transfer_count[0][11] ),
    .A3(_0589_),
    .B1(_0584_),
    .Y(_0597_));
 sky130_fd_sc_hd__o21ai_0 _2290_ (.A1(_0558_),
    .A2(_0597_),
    .B1(\transfer_count[0][13] ),
    .Y(_0598_));
 sky130_fd_sc_hd__o31ai_1 _2291_ (.A1(\transfer_count[0][13] ),
    .A2(_0995_),
    .A3(_0556_),
    .B1(_0598_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand3_1 _2292_ (.A(_1006_),
    .B(_1007_),
    .C(_0581_),
    .Y(_0599_));
 sky130_fd_sc_hd__xor2_1 _2293_ (.A(\transfer_count[0][14] ),
    .B(_0599_),
    .X(_1234_));
 sky130_fd_sc_hd__nand2_1 _2294_ (.A(\transfer_count[0][14] ),
    .B(_0558_),
    .Y(_0600_));
 sky130_fd_sc_hd__o21ai_0 _2295_ (.A1(_0556_),
    .A2(_1234_),
    .B1(_0600_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _2296_ (.A(_1015_),
    .B(_0149_),
    .Y(_0601_));
 sky130_fd_sc_hd__o21ai_0 _2297_ (.A1(_1015_),
    .A2(_0584_),
    .B1(_0592_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _2298_ (.A(\transfer_count[0][15] ),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__o21ai_0 _2299_ (.A1(\transfer_count[0][15] ),
    .A2(_0601_),
    .B1(_0603_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_2 _2300_ (.A(_1008_),
    .B(_0580_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_1 _2301_ (.A(_0150_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__o21ai_0 _2302_ (.A1(_0555_),
    .A2(_0604_),
    .B1(_0592_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _2303_ (.A(_1003_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__o21ai_0 _2304_ (.A1(_1003_),
    .A2(_0605_),
    .B1(_0607_),
    .Y(_0020_));
 sky130_fd_sc_hd__a31oi_1 _2305_ (.A1(\transfer_count[0][15] ),
    .A2(_1003_),
    .A3(_1015_),
    .B1(_0584_),
    .Y(_0608_));
 sky130_fd_sc_hd__o21ai_0 _2306_ (.A1(_0563_),
    .A2(_0608_),
    .B1(\transfer_count[0][17] ),
    .Y(_0609_));
 sky130_fd_sc_hd__o31ai_1 _2307_ (.A1(\transfer_count[0][17] ),
    .A2(_0146_),
    .A3(_0556_),
    .B1(_0609_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand3_1 _2308_ (.A(\transfer_count[0][17] ),
    .B(_1003_),
    .C(_0604_),
    .Y(_0610_));
 sky130_fd_sc_hd__a31oi_1 _2309_ (.A1(\transfer_count[0][17] ),
    .A2(_1003_),
    .A3(_0604_),
    .B1(_0584_),
    .Y(_0611_));
 sky130_fd_sc_hd__o21ai_0 _2310_ (.A1(_0563_),
    .A2(_0611_),
    .B1(\transfer_count[0][18] ),
    .Y(_0612_));
 sky130_fd_sc_hd__o31ai_1 _2311_ (.A1(\transfer_count[0][18] ),
    .A2(_0560_),
    .A3(_0610_),
    .B1(_0612_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand3_1 _2312_ (.A(\transfer_count[0][18] ),
    .B(\transfer_count[0][17] ),
    .C(_1003_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor3_1 _2313_ (.A(_0993_),
    .B(_0613_),
    .C(_1008_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _2314_ (.A(_0150_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__o21ai_0 _2315_ (.A1(_0555_),
    .A2(_0614_),
    .B1(_0592_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _2316_ (.A(\transfer_count[0][19] ),
    .B(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__o21ai_0 _2317_ (.A1(\transfer_count[0][19] ),
    .A2(_0615_),
    .B1(_0617_),
    .Y(_0023_));
 sky130_fd_sc_hd__nand3_1 _2318_ (.A(\transfer_count[0][19] ),
    .B(_1004_),
    .C(_0604_),
    .Y(_0618_));
 sky130_fd_sc_hd__a31oi_1 _2319_ (.A1(\transfer_count[0][19] ),
    .A2(_1004_),
    .A3(_0604_),
    .B1(_0584_),
    .Y(_0619_));
 sky130_fd_sc_hd__o21ai_0 _2320_ (.A1(_0563_),
    .A2(_0619_),
    .B1(\transfer_count[0][20] ),
    .Y(_0620_));
 sky130_fd_sc_hd__o31ai_1 _2321_ (.A1(\transfer_count[0][20] ),
    .A2(_0560_),
    .A3(_0618_),
    .B1(_0620_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2b_1 _2322_ (.A_N(_1016_),
    .B(_0149_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21oi_1 _2323_ (.A1(_1016_),
    .A2(_0149_),
    .B1(\transfer_count[0][21] ),
    .Y(_0622_));
 sky130_fd_sc_hd__a31oi_1 _2324_ (.A1(\transfer_count[0][21] ),
    .A2(_0592_),
    .A3(_0621_),
    .B1(_0622_),
    .Y(_0026_));
 sky130_fd_sc_hd__nor3_4 _2325_ (.A(_1005_),
    .B(_1008_),
    .C(_0580_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _2326_ (.A(_0150_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nor2_1 _2327_ (.A(_0584_),
    .B(_0623_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21ai_0 _2328_ (.A1(_0557_),
    .A2(_0625_),
    .B1(_0999_),
    .Y(_0626_));
 sky130_fd_sc_hd__o21ai_0 _2329_ (.A1(_0999_),
    .A2(_0624_),
    .B1(_0626_),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _2330_ (.A(_0999_),
    .B(_1009_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _2331_ (.A(_0149_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__a31oi_1 _2332_ (.A1(_0999_),
    .A2(_1009_),
    .A3(_0149_),
    .B1(\transfer_count[0][23] ),
    .Y(_0629_));
 sky130_fd_sc_hd__a31oi_1 _2333_ (.A1(\transfer_count[0][23] ),
    .A2(_0592_),
    .A3(_0628_),
    .B1(_0629_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand3_1 _2334_ (.A(\transfer_count[0][23] ),
    .B(_0999_),
    .C(_0623_),
    .Y(_0630_));
 sky130_fd_sc_hd__a31oi_1 _2335_ (.A1(\transfer_count[0][23] ),
    .A2(_0999_),
    .A3(_0623_),
    .B1(_0584_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21ai_0 _2336_ (.A1(_0563_),
    .A2(_0631_),
    .B1(\transfer_count[0][24] ),
    .Y(_0632_));
 sky130_fd_sc_hd__o31ai_1 _2337_ (.A1(\transfer_count[0][24] ),
    .A2(_0560_),
    .A3(_0630_),
    .B1(_0632_),
    .Y(_0029_));
 sky130_fd_sc_hd__a21oi_1 _2338_ (.A1(_1011_),
    .A2(_1009_),
    .B1(_0564_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ai_0 _2339_ (.A1(_0563_),
    .A2(_0633_),
    .B1(\transfer_count[0][25] ),
    .Y(_0634_));
 sky130_fd_sc_hd__o31ai_1 _2340_ (.A1(\transfer_count[0][25] ),
    .A2(_1012_),
    .A3(_0560_),
    .B1(_0634_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _2341_ (.A(_1001_),
    .B(_0623_),
    .Y(_0635_));
 sky130_fd_sc_hd__a21oi_1 _2342_ (.A1(_1001_),
    .A2(_0623_),
    .B1(_0564_),
    .Y(_0636_));
 sky130_fd_sc_hd__o21ai_0 _2343_ (.A1(_0563_),
    .A2(_0636_),
    .B1(\transfer_count[0][26] ),
    .Y(_0637_));
 sky130_fd_sc_hd__o31ai_1 _2344_ (.A1(\transfer_count[0][26] ),
    .A2(_0560_),
    .A3(_0635_),
    .B1(_0637_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand3_1 _2345_ (.A(\transfer_count[0][26] ),
    .B(_1001_),
    .C(_1009_),
    .Y(_0638_));
 sky130_fd_sc_hd__a31oi_1 _2346_ (.A1(\transfer_count[0][26] ),
    .A2(_1001_),
    .A3(_1009_),
    .B1(_0584_),
    .Y(_0639_));
 sky130_fd_sc_hd__o21ai_0 _2347_ (.A1(_0563_),
    .A2(_0639_),
    .B1(\transfer_count[0][27] ),
    .Y(_0640_));
 sky130_fd_sc_hd__o31ai_1 _2348_ (.A1(\transfer_count[0][27] ),
    .A2(_0560_),
    .A3(_0638_),
    .B1(_0640_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand3_1 _2349_ (.A(\transfer_count[0][27] ),
    .B(\transfer_count[0][26] ),
    .C(_1001_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor4_1 _2350_ (.A(_0641_),
    .B(_1005_),
    .C(_1008_),
    .D(_0580_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_1 _2351_ (.A(_0150_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__o21ai_0 _2352_ (.A1(_0555_),
    .A2(_0642_),
    .B1(_0592_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _2353_ (.A(\transfer_count[0][28] ),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ai_0 _2354_ (.A1(\transfer_count[0][28] ),
    .A2(_0643_),
    .B1(_0645_),
    .Y(_0033_));
 sky130_fd_sc_hd__nand2_1 _2355_ (.A(_1010_),
    .B(_0149_),
    .Y(_0646_));
 sky130_fd_sc_hd__a31oi_1 _2356_ (.A1(_1002_),
    .A2(_1009_),
    .A3(_0149_),
    .B1(\transfer_count[0][29] ),
    .Y(_0647_));
 sky130_fd_sc_hd__a31oi_1 _2357_ (.A1(\transfer_count[0][29] ),
    .A2(_0592_),
    .A3(_0646_),
    .B1(_0647_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand3_1 _2358_ (.A(\transfer_count[0][29] ),
    .B(_1002_),
    .C(_0623_),
    .Y(_0648_));
 sky130_fd_sc_hd__a31oi_1 _2359_ (.A1(\transfer_count[0][29] ),
    .A2(_1002_),
    .A3(_0623_),
    .B1(_0584_),
    .Y(_0649_));
 sky130_fd_sc_hd__o21ai_0 _2360_ (.A1(_0563_),
    .A2(_0649_),
    .B1(\transfer_count[0][30] ),
    .Y(_0650_));
 sky130_fd_sc_hd__o31ai_1 _2361_ (.A1(\transfer_count[0][30] ),
    .A2(_0564_),
    .A3(_0648_),
    .B1(_0650_),
    .Y(_0036_));
 sky130_fd_sc_hd__and3_1 _2362_ (.A(\transfer_count[0][30] ),
    .B(\transfer_count[0][29] ),
    .C(_1002_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _2363_ (.A(_1009_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__a21oi_1 _2364_ (.A1(_1009_),
    .A2(_0651_),
    .B1(_0564_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21ai_0 _2365_ (.A1(_0563_),
    .A2(_0653_),
    .B1(\transfer_count[0][31] ),
    .Y(_0654_));
 sky130_fd_sc_hd__o31ai_1 _2366_ (.A1(\transfer_count[0][31] ),
    .A2(_0564_),
    .A3(_0652_),
    .B1(_0654_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_1 _2367_ (.A(\active_channel_count[0] ),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2b_1 _2368_ (.A_N(_0980_),
    .B(_0981_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2b_2 _2369_ (.A_N(_0981_),
    .B(_0980_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _2370_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(net2),
    .B(net146),
    .Y(_0658_));
 sky130_fd_sc_hd__a21oi_1 _2372_ (.A1(\channel_state[0][2] ),
    .A2(_0657_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nor2b_1 _2373_ (.A(_0825_),
    .B_N(_0826_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2b_1 _2374_ (.A_N(\channel_state[1][1] ),
    .B(\channel_state[1][0] ),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2b_1 _2375_ (.A_N(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _2376_ (.A(net147),
    .B(net3),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _2377_ (.A1(_0445_),
    .A2(_0662_),
    .B1(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__inv_1 _2378_ (.A(\channel_state[3][1] ),
    .Y(_0665_));
 sky130_fd_sc_hd__nor2_1 _2379_ (.A(\channel_state[3][0] ),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _2380_ (.A(_0976_),
    .B(_0665_),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2b_1 _2381_ (.A_N(_0666_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(net149),
    .B(net5),
    .Y(_0669_));
 sky130_fd_sc_hd__a21oi_4 _2383_ (.A1(_0920_),
    .A2(_0668_),
    .B1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__clkbuf_2 _2384_ (.A(\channel_state[2][1] ),
    .X(_0671_));
 sky130_fd_sc_hd__nor2b_1 _2385_ (.A(\channel_state[2][0] ),
    .B_N(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2b_1 _2386_ (.A_N(\channel_state[2][1] ),
    .B(\channel_state[2][0] ),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2b_1 _2387_ (.A_N(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _2388_ (.A(net148),
    .B(net4),
    .Y(_0675_));
 sky130_fd_sc_hd__a21oi_1 _2389_ (.A1(_0308_),
    .A2(_0674_),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor4_2 _2390_ (.A(_0659_),
    .B(_0664_),
    .C(_0670_),
    .D(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nor2_1 _2391_ (.A(\active_channel_count[0] ),
    .B(_0677_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2b_1 _2392_ (.A(_0677_),
    .B_N(_1306_),
    .Y(_0001_));
 sky130_fd_sc_hd__xnor2_1 _2393_ (.A(_1307_),
    .B(\active_channel_count[2] ),
    .Y(_0678_));
 sky130_fd_sc_hd__nor2_1 _2394_ (.A(_0677_),
    .B(_0678_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand3_1 _2395_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[2] ),
    .C(\active_channel_count[1] ),
    .Y(_0679_));
 sky130_fd_sc_hd__xor2_1 _2396_ (.A(\active_channel_count[3] ),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _2397_ (.A(_0677_),
    .B(_0680_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _2398_ (.A(net134),
    .B(_0553_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2b_1 _2399_ (.A_N(_0553_),
    .B(net142),
    .Y(_0682_));
 sky130_fd_sc_hd__o221ai_1 _2400_ (.A1(_0656_),
    .A2(_0681_),
    .B1(_0682_),
    .B2(_0655_),
    .C1(_0558_),
    .Y(_1030_));
 sky130_fd_sc_hd__nor2_2 _2401_ (.A(_0553_),
    .B(_0656_),
    .Y(_1019_));
 sky130_fd_sc_hd__o22ai_1 _2402_ (.A1(_0982_),
    .A2(_0655_),
    .B1(_0656_),
    .B2(_0553_),
    .Y(_1031_));
 sky130_fd_sc_hd__a21o_1 _2403_ (.A1(net134),
    .A2(_0657_),
    .B1(_0147_),
    .X(_0683_));
 sky130_fd_sc_hd__nand2_1 _2404_ (.A(_0980_),
    .B(_0981_),
    .Y(_0684_));
 sky130_fd_sc_hd__o211ai_1 _2405_ (.A1(net134),
    .A2(_0554_),
    .B1(_0684_),
    .C1(_0553_),
    .Y(_0685_));
 sky130_fd_sc_hd__o21ai_0 _2406_ (.A1(_0553_),
    .A2(_0684_),
    .B1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__o21a_1 _2407_ (.A1(_0201_),
    .A2(_0683_),
    .B1(_0686_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2b_1 _2408_ (.A_N(_0826_),
    .B(net135),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _2409_ (.A(_0445_),
    .B(_0825_),
    .Y(_0688_));
 sky130_fd_sc_hd__inv_1 _2410_ (.A(_0445_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand3_1 _2411_ (.A(_0689_),
    .B(net143),
    .C(_0660_),
    .Y(_0690_));
 sky130_fd_sc_hd__o211ai_1 _2412_ (.A1(_0687_),
    .A2(_0688_),
    .B1(_0690_),
    .C1(_0455_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_2 _2413_ (.A(_0445_),
    .B(_0661_),
    .Y(_1018_));
 sky130_fd_sc_hd__a22o_1 _2414_ (.A1(net135),
    .A2(_0660_),
    .B1(_0662_),
    .B2(_0689_),
    .X(_1028_));
 sky130_fd_sc_hd__inv_1 _2415_ (.A(net139),
    .Y(_0691_));
 sky130_fd_sc_hd__a311oi_1 _2416_ (.A1(_0445_),
    .A2(_0825_),
    .A3(net135),
    .B1(_0826_),
    .C1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2b_1 _2417_ (.A(net135),
    .B_N(_0826_),
    .Y(_0693_));
 sky130_fd_sc_hd__o21ai_0 _2418_ (.A1(_0825_),
    .A2(_0693_),
    .B1(_0687_),
    .Y(_0694_));
 sky130_fd_sc_hd__and3_1 _2419_ (.A(_0689_),
    .B(_0825_),
    .C(_0826_),
    .X(_0695_));
 sky130_fd_sc_hd__a21oi_1 _2420_ (.A1(_0445_),
    .A2(_0694_),
    .B1(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a21oi_1 _2421_ (.A1(_0880_),
    .A2(_0692_),
    .B1(_0696_),
    .Y(_1029_));
 sky130_fd_sc_hd__nand2b_1 _2422_ (.A_N(_0671_),
    .B(net136),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _2423_ (.A(_0308_),
    .B(\channel_state[2][0] ),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_1 _2424_ (.A(net144),
    .B(_0672_),
    .Y(_0699_));
 sky130_fd_sc_hd__o221ai_1 _2425_ (.A1(_0697_),
    .A2(_0698_),
    .B1(_0699_),
    .B2(_0308_),
    .C1(_0313_),
    .Y(_1024_));
 sky130_fd_sc_hd__nor2_2 _2426_ (.A(_0308_),
    .B(_0673_),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_1 _2427_ (.A(_0308_),
    .Y(_0700_));
 sky130_fd_sc_hd__a22o_1 _2428_ (.A1(net136),
    .A2(_0672_),
    .B1(_0674_),
    .B2(_0700_),
    .X(_1025_));
 sky130_fd_sc_hd__nand3_1 _2429_ (.A(_0700_),
    .B(\channel_state[2][0] ),
    .C(_0671_),
    .Y(_0701_));
 sky130_fd_sc_hd__nor2b_1 _2430_ (.A(net136),
    .B_N(_0671_),
    .Y(_0702_));
 sky130_fd_sc_hd__o21ai_0 _2431_ (.A1(\channel_state[2][0] ),
    .A2(_0702_),
    .B1(_0697_),
    .Y(_0703_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(_0308_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand2_1 _2433_ (.A(_0701_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__and3_1 _2434_ (.A(_1311_),
    .B(_1314_),
    .C(_1317_),
    .X(_0706_));
 sky130_fd_sc_hd__a211oi_1 _2435_ (.A1(_1331_),
    .A2(_1329_),
    .B1(_1325_),
    .C1(_1328_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21ai_0 _2436_ (.A1(_1326_),
    .A2(_1325_),
    .B1(_1323_),
    .Y(_0708_));
 sky130_fd_sc_hd__nor2_1 _2437_ (.A(_1319_),
    .B(_1322_),
    .Y(_0709_));
 sky130_fd_sc_hd__o21ai_0 _2438_ (.A1(_0707_),
    .A2(_0708_),
    .B1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o211ai_1 _2439_ (.A1(_1319_),
    .A2(_1320_),
    .B1(_0706_),
    .C1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21oi_1 _2440_ (.A1(_1314_),
    .A2(_1316_),
    .B1(_1313_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2b_1 _2441_ (.A(_0712_),
    .B_N(_1311_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21oi_1 _2442_ (.A1(_1335_),
    .A2(_1337_),
    .B1(_1334_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand4_2 _2443_ (.A(_1320_),
    .B(_1326_),
    .C(_1332_),
    .D(_1329_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand4_2 _2444_ (.A(_1311_),
    .B(_1323_),
    .C(_1314_),
    .D(_1317_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor3_1 _2445_ (.A(_0714_),
    .B(_0715_),
    .C(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor3_1 _2446_ (.A(_1310_),
    .B(_0713_),
    .C(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21oi_1 _2447_ (.A1(_1355_),
    .A2(_1353_),
    .B1(_1352_),
    .Y(_0719_));
 sky130_fd_sc_hd__nand3_1 _2448_ (.A(_1347_),
    .B(_1344_),
    .C(_1350_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand3_1 _2449_ (.A(_1347_),
    .B(_1344_),
    .C(_1349_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _2450_ (.A(_1344_),
    .B(_1346_),
    .Y(_0722_));
 sky130_fd_sc_hd__o211ai_1 _2451_ (.A1(_0719_),
    .A2(_0720_),
    .B1(_0721_),
    .C1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand2_1 _2452_ (.A(_1335_),
    .B(_1338_),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _2453_ (.A(_1341_),
    .B(_1340_),
    .Y(_0725_));
 sky130_fd_sc_hd__nor4_1 _2454_ (.A(_0715_),
    .B(_0716_),
    .C(_0724_),
    .D(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o31ai_1 _2455_ (.A1(_1343_),
    .A2(_1340_),
    .A3(_0723_),
    .B1(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__and3_1 _2456_ (.A(_0711_),
    .B(_0718_),
    .C(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2b_1 _2457_ (.A(_1406_),
    .B_N(_1403_),
    .Y(_0729_));
 sky130_fd_sc_hd__o211ai_1 _2458_ (.A1(_1402_),
    .A2(_0729_),
    .B1(_1395_),
    .C1(_1398_),
    .Y(_0730_));
 sky130_fd_sc_hd__a21oi_1 _2459_ (.A1(_1395_),
    .A2(_1397_),
    .B1(_1394_),
    .Y(_0731_));
 sky130_fd_sc_hd__nand4_1 _2460_ (.A(_1383_),
    .B(_1386_),
    .C(_1392_),
    .D(_1389_),
    .Y(_0732_));
 sky130_fd_sc_hd__a21oi_1 _2461_ (.A1(_0730_),
    .A2(_0731_),
    .B1(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _2462_ (.A(_1383_),
    .B(_1386_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _2463_ (.A1(_1391_),
    .A2(_1389_),
    .B1(_1388_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2464_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a21oi_1 _2465_ (.A1(_1359_),
    .A2(_1361_),
    .B1(_1358_),
    .Y(_0737_));
 sky130_fd_sc_hd__a21oi_1 _2466_ (.A1(_1383_),
    .A2(_1385_),
    .B1(_1382_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _2467_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand4_1 _2468_ (.A(_1368_),
    .B(_1374_),
    .C(_1380_),
    .D(_1365_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand4_1 _2469_ (.A(_1359_),
    .B(_1371_),
    .C(_1362_),
    .D(_1377_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21ai_0 _2470_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0737_),
    .Y(_0742_));
 sky130_fd_sc_hd__and4_1 _2471_ (.A(_1347_),
    .B(_1344_),
    .C(_1356_),
    .D(_1341_),
    .X(_0743_));
 sky130_fd_sc_hd__nand3_1 _2472_ (.A(_1350_),
    .B(_1353_),
    .C(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor4_2 _2473_ (.A(_0715_),
    .B(_0716_),
    .C(_0724_),
    .D(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__o311ai_2 _2474_ (.A1(_0733_),
    .A2(_0736_),
    .A3(_0739_),
    .B1(_0742_),
    .C1(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__a21o_1 _2475_ (.A1(_1379_),
    .A2(_1377_),
    .B1(_1376_),
    .X(_0747_));
 sky130_fd_sc_hd__a21oi_1 _2476_ (.A1(_1374_),
    .A2(_0747_),
    .B1(_1373_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _2477_ (.A(_1371_),
    .B(_1368_),
    .Y(_0749_));
 sky130_fd_sc_hd__a211oi_1 _2478_ (.A1(_1368_),
    .A2(_1370_),
    .B1(_1364_),
    .C1(_1367_),
    .Y(_0750_));
 sky130_fd_sc_hd__o21ai_0 _2479_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__o211a_1 _2480_ (.A1(_1365_),
    .A2(_1364_),
    .B1(_1359_),
    .C1(_1362_),
    .X(_0752_));
 sky130_fd_sc_hd__nand3_1 _2481_ (.A(_0751_),
    .B(_0752_),
    .C(_0745_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand4_1 _2482_ (.A(_0705_),
    .B(_0728_),
    .C(_0746_),
    .D(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand4_1 _2483_ (.A(_1395_),
    .B(_1403_),
    .C(_1407_),
    .D(_1398_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor4_1 _2484_ (.A(_0732_),
    .B(_0740_),
    .C(_0741_),
    .D(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _2485_ (.A(net140),
    .B(_0671_),
    .Y(_0757_));
 sky130_fd_sc_hd__a21oi_1 _2486_ (.A1(net136),
    .A2(_0671_),
    .B1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2b_1 _2487_ (.A(_0671_),
    .B_N(net136),
    .Y(_0759_));
 sky130_fd_sc_hd__mux2i_1 _2488_ (.A0(_0671_),
    .A1(_0759_),
    .S(_0308_),
    .Y(_0760_));
 sky130_fd_sc_hd__o22ai_1 _2489_ (.A1(_0301_),
    .A2(_0758_),
    .B1(_0760_),
    .B2(_0307_),
    .Y(_0761_));
 sky130_fd_sc_hd__a31oi_1 _2490_ (.A1(_0705_),
    .A2(_0745_),
    .A3(_0756_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _2491_ (.A(_0754_),
    .B(_0762_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _2492_ (.A(_0920_),
    .B(_0667_),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _2493_ (.A(net137),
    .B(_0665_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _2494_ (.A(_0920_),
    .B(_0976_),
    .Y(_0764_));
 sky130_fd_sc_hd__inv_1 _2495_ (.A(_0920_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand3_1 _2496_ (.A(_0765_),
    .B(net145),
    .C(_0666_),
    .Y(_0766_));
 sky130_fd_sc_hd__o211ai_1 _2497_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0766_),
    .C1(_0208_),
    .Y(_1021_));
 sky130_fd_sc_hd__a22o_1 _2498_ (.A1(net137),
    .A2(_0666_),
    .B1(_0668_),
    .B2(_0765_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _2499_ (.A(net137),
    .B(_0665_),
    .Y(_0767_));
 sky130_fd_sc_hd__o21ai_0 _2500_ (.A1(_0976_),
    .A2(_0767_),
    .B1(_0763_),
    .Y(_0768_));
 sky130_fd_sc_hd__and3_1 _2501_ (.A(_0765_),
    .B(_0976_),
    .C(\channel_state[3][1] ),
    .X(_0769_));
 sky130_fd_sc_hd__a21oi_1 _2502_ (.A1(_0920_),
    .A2(_0768_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__nor2b_1 _2503_ (.A(\channel_state[3][1] ),
    .B_N(net137),
    .Y(_0771_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(\channel_state[3][1] ),
    .A1(_0771_),
    .S(_0920_),
    .X(_0772_));
 sky130_fd_sc_hd__a2111oi_0 _2505_ (.A1(net141),
    .A2(_0665_),
    .B1(_0767_),
    .C1(_0765_),
    .D1(_0976_),
    .Y(_0773_));
 sky130_fd_sc_hd__a21oi_1 _2506_ (.A1(_0976_),
    .A2(_0772_),
    .B1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__o31ai_1 _2507_ (.A1(_0954_),
    .A2(_0975_),
    .A3(_0770_),
    .B1(_0774_),
    .Y(_1023_));
 sky130_fd_sc_hd__o21a_1 _2508_ (.A1(net142),
    .A2(_0655_),
    .B1(_0656_),
    .X(_0775_));
 sky130_fd_sc_hd__nor2_2 _2509_ (.A(_0553_),
    .B(_0775_),
    .Y(_1442_));
 sky130_fd_sc_hd__nor2_1 _2510_ (.A(_0980_),
    .B(_0983_),
    .Y(_0776_));
 sky130_fd_sc_hd__a21oi_1 _2511_ (.A1(_0980_),
    .A2(_0982_),
    .B1(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__o21ai_0 _2512_ (.A1(_0981_),
    .A2(_0777_),
    .B1(net150),
    .Y(_0778_));
 sky130_fd_sc_hd__a21bo_1 _2513_ (.A1(_0150_),
    .A2(_0201_),
    .B1_N(_0778_),
    .X(_1441_));
 sky130_fd_sc_hd__nand2b_1 _2514_ (.A_N(net143),
    .B(_0660_),
    .Y(_0779_));
 sky130_fd_sc_hd__a21oi_2 _2515_ (.A1(_0661_),
    .A2(_0779_),
    .B1(_0445_),
    .Y(_1440_));
 sky130_fd_sc_hd__o22a_1 _2516_ (.A1(_0825_),
    .A2(_0882_),
    .B1(_0688_),
    .B2(net135),
    .X(_0780_));
 sky130_fd_sc_hd__o21ai_0 _2517_ (.A1(_0826_),
    .A2(_0780_),
    .B1(net151),
    .Y(_0781_));
 sky130_fd_sc_hd__o21ai_0 _2518_ (.A1(_0452_),
    .A2(_0880_),
    .B1(_0781_),
    .Y(_1439_));
 sky130_fd_sc_hd__o22a_1 _2519_ (.A1(_0976_),
    .A2(_0978_),
    .B1(_0764_),
    .B2(net137),
    .X(_0782_));
 sky130_fd_sc_hd__o21ai_0 _2520_ (.A1(\channel_state[3][1] ),
    .A2(_0782_),
    .B1(net153),
    .Y(_0783_));
 sky130_fd_sc_hd__o31ai_1 _2521_ (.A1(_0223_),
    .A2(_0954_),
    .A3(_0975_),
    .B1(_0783_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2b_1 _2522_ (.A_N(net144),
    .B(_0672_),
    .Y(_0784_));
 sky130_fd_sc_hd__a21oi_2 _2523_ (.A1(_0673_),
    .A2(_0784_),
    .B1(_0308_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand4_1 _2524_ (.A(_0306_),
    .B(_0728_),
    .C(_0746_),
    .D(_0753_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand3_1 _2525_ (.A(_0316_),
    .B(_0745_),
    .C(_0756_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21ba_1 _2526_ (.A1(net136),
    .A2(_0698_),
    .B1_N(_0310_),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_0 _2527_ (.A1(_0671_),
    .A2(_0787_),
    .B1(net152),
    .Y(_0788_));
 sky130_fd_sc_hd__nand3_1 _2528_ (.A(_0785_),
    .B(_0786_),
    .C(_0788_),
    .Y(_1436_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(\active_channel_count[2] ),
    .B(\active_channel_count[3] ),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _2530_ (.A(_1305_),
    .B(_0789_),
    .Y(_0012_));
 sky130_fd_sc_hd__a22oi_1 _2531_ (.A1(_0977_),
    .A2(_0771_),
    .B1(_0767_),
    .B2(_0920_),
    .Y(_0790_));
 sky130_fd_sc_hd__o21a_1 _2532_ (.A1(_0976_),
    .A2(_0790_),
    .B1(net157),
    .X(_0011_));
 sky130_fd_sc_hd__a22oi_1 _2533_ (.A1(_0309_),
    .A2(_0759_),
    .B1(_0702_),
    .B2(_0308_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21a_1 _2534_ (.A1(\channel_state[2][0] ),
    .A2(_0791_),
    .B1(net156),
    .X(_0010_));
 sky130_fd_sc_hd__o211a_1 _2535_ (.A1(net148),
    .A2(_0311_),
    .B1(_0785_),
    .C1(_0786_),
    .X(_0006_));
 sky130_fd_sc_hd__nor2b_1 _2536_ (.A(_0826_),
    .B_N(net135),
    .Y(_0792_));
 sky130_fd_sc_hd__a22oi_1 _2537_ (.A1(_0881_),
    .A2(_0792_),
    .B1(_0693_),
    .B2(_0445_),
    .Y(_0793_));
 sky130_fd_sc_hd__o21a_1 _2538_ (.A1(_0825_),
    .A2(_0793_),
    .B1(net155),
    .X(_0009_));
 sky130_fd_sc_hd__inv_1 _2539_ (.A(net129),
    .Y(_1200_));
 sky130_fd_sc_hd__inv_1 _2540_ (.A(net6),
    .Y(_1204_));
 sky130_fd_sc_hd__xnor2_1 _2541_ (.A(\transfer_count[2][30] ),
    .B(_0438_),
    .Y(_1312_));
 sky130_fd_sc_hd__xor2_1 _2542_ (.A(\transfer_count[2][26] ),
    .B(_0423_),
    .X(_1324_));
 sky130_fd_sc_hd__inv_1 _2543_ (.A(net94),
    .Y(_1404_));
 sky130_fd_sc_hd__inv_1 _2544_ (.A(net59),
    .Y(_1408_));
 sky130_fd_sc_hd__xnor2_1 _2545_ (.A(\transfer_count[1][8] ),
    .B(_0477_),
    .Y(_1054_));
 sky130_fd_sc_hd__nor2_1 _2546_ (.A(_0820_),
    .B(_0549_),
    .Y(_0794_));
 sky130_fd_sc_hd__xnor2_1 _2547_ (.A(\transfer_count[1][31] ),
    .B(_0794_),
    .Y(_1057_));
 sky130_fd_sc_hd__xor2_1 _2548_ (.A(\transfer_count[1][30] ),
    .B(_0545_),
    .X(_1060_));
 sky130_fd_sc_hd__xnor2_1 _2549_ (.A(\transfer_count[1][28] ),
    .B(_0540_),
    .Y(_1066_));
 sky130_fd_sc_hd__xnor2_1 _2550_ (.A(_0534_),
    .B(_0535_),
    .Y(_1069_));
 sky130_fd_sc_hd__xor2_1 _2551_ (.A(\transfer_count[1][26] ),
    .B(_0530_),
    .X(_1072_));
 sky130_fd_sc_hd__xor2_1 _2552_ (.A(\transfer_count[1][24] ),
    .B(_0525_),
    .X(_1078_));
 sky130_fd_sc_hd__xor2_1 _2553_ (.A(\transfer_count[1][23] ),
    .B(_0522_),
    .X(_1081_));
 sky130_fd_sc_hd__xor2_1 _2554_ (.A(\transfer_count[1][22] ),
    .B(_0519_),
    .X(_1084_));
 sky130_fd_sc_hd__xor2_1 _2555_ (.A(\transfer_count[1][20] ),
    .B(_0513_),
    .X(_1090_));
 sky130_fd_sc_hd__xnor2_1 _2556_ (.A(\transfer_count[1][19] ),
    .B(_0510_),
    .Y(_1093_));
 sky130_fd_sc_hd__xor2_1 _2557_ (.A(\transfer_count[1][18] ),
    .B(_0504_),
    .X(_1096_));
 sky130_fd_sc_hd__xnor2_1 _2558_ (.A(\transfer_count[1][16] ),
    .B(_0496_),
    .Y(_1102_));
 sky130_fd_sc_hd__xnor2_1 _2559_ (.A(\transfer_count[3][31] ),
    .B(_0299_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_1 _2560_ (.A(\transfer_count[3][30] ),
    .B(_0295_),
    .Y(_1108_));
 sky130_fd_sc_hd__xnor2_1 _2561_ (.A(\transfer_count[3][28] ),
    .B(_0288_),
    .Y(_1114_));
 sky130_fd_sc_hd__xnor2_1 _2562_ (.A(\transfer_count[3][26] ),
    .B(_0281_),
    .Y(_1120_));
 sky130_fd_sc_hd__xor2_1 _2563_ (.A(_0884_),
    .B(_0274_),
    .X(_1126_));
 sky130_fd_sc_hd__xnor2_1 _2564_ (.A(\transfer_count[3][22] ),
    .B(_0268_),
    .Y(_1132_));
 sky130_fd_sc_hd__xnor2_1 _2565_ (.A(\transfer_count[3][20] ),
    .B(_0263_),
    .Y(_1138_));
 sky130_fd_sc_hd__xor2_1 _2566_ (.A(\transfer_count[3][18] ),
    .B(_0259_),
    .X(_1144_));
 sky130_fd_sc_hd__xor2_1 _2567_ (.A(\transfer_count[3][17] ),
    .B(_0256_),
    .X(_1147_));
 sky130_fd_sc_hd__xnor2_1 _2568_ (.A(\transfer_count[3][16] ),
    .B(_0252_),
    .Y(_1150_));
 sky130_fd_sc_hd__xnor2_1 _2569_ (.A(\transfer_count[3][14] ),
    .B(_0246_),
    .Y(_1156_));
 sky130_fd_sc_hd__xor2_1 _2570_ (.A(\transfer_count[3][6] ),
    .B(_0225_),
    .X(_1180_));
 sky130_fd_sc_hd__xnor2_1 _2571_ (.A(\transfer_count[3][2] ),
    .B(_0211_),
    .Y(_1192_));
 sky130_fd_sc_hd__xnor2_1 _2572_ (.A(\transfer_count[0][3] ),
    .B(_0987_),
    .Y(_1213_));
 sky130_fd_sc_hd__xnor2_1 _2573_ (.A(\transfer_count[0][2] ),
    .B(_1208_),
    .Y(_1216_));
 sky130_fd_sc_hd__xnor2_1 _2574_ (.A(_0991_),
    .B(_0997_),
    .Y(_1219_));
 sky130_fd_sc_hd__xor2_1 _2575_ (.A(\transfer_count[0][6] ),
    .B(_0573_),
    .X(_1222_));
 sky130_fd_sc_hd__xnor2_1 _2576_ (.A(\transfer_count[0][15] ),
    .B(_1015_),
    .Y(_1231_));
 sky130_fd_sc_hd__xnor2_1 _2577_ (.A(\transfer_count[0][11] ),
    .B(_0589_),
    .Y(_1243_));
 sky130_fd_sc_hd__xor2_1 _2578_ (.A(_0989_),
    .B(_0580_),
    .X(_1252_));
 sky130_fd_sc_hd__xor2_1 _2579_ (.A(\transfer_count[0][31] ),
    .B(_0652_),
    .X(_1255_));
 sky130_fd_sc_hd__xor2_1 _2580_ (.A(\transfer_count[0][30] ),
    .B(_0648_),
    .X(_1258_));
 sky130_fd_sc_hd__xnor2_1 _2581_ (.A(\transfer_count[0][28] ),
    .B(_0642_),
    .Y(_1264_));
 sky130_fd_sc_hd__xor2_1 _2582_ (.A(\transfer_count[0][27] ),
    .B(_0638_),
    .X(_1267_));
 sky130_fd_sc_hd__xor2_1 _2583_ (.A(\transfer_count[0][26] ),
    .B(_0635_),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _2584_ (.A(\transfer_count[0][24] ),
    .B(_0630_),
    .X(_1276_));
 sky130_fd_sc_hd__xor2_1 _2585_ (.A(\transfer_count[0][23] ),
    .B(_0627_),
    .X(_1279_));
 sky130_fd_sc_hd__xnor2_1 _2586_ (.A(_0999_),
    .B(_0623_),
    .Y(_1282_));
 sky130_fd_sc_hd__xor2_1 _2587_ (.A(\transfer_count[0][20] ),
    .B(_0618_),
    .X(_1288_));
 sky130_fd_sc_hd__xnor2_1 _2588_ (.A(\transfer_count[0][19] ),
    .B(_0614_),
    .Y(_1291_));
 sky130_fd_sc_hd__xor2_1 _2589_ (.A(\transfer_count[0][18] ),
    .B(_0610_),
    .X(_1294_));
 sky130_fd_sc_hd__xnor2_1 _2590_ (.A(_1003_),
    .B(_0604_),
    .Y(_1300_));
 sky130_fd_sc_hd__inv_1 _2591_ (.A(\active_channel_count[1] ),
    .Y(_1304_));
 sky130_fd_sc_hd__xor2_1 _2592_ (.A(\transfer_count[2][31] ),
    .B(_0442_),
    .X(_1309_));
 sky130_fd_sc_hd__xor2_1 _2593_ (.A(\transfer_count[2][28] ),
    .B(_0431_),
    .X(_1318_));
 sky130_fd_sc_hd__xor2_1 _2594_ (.A(\transfer_count[2][24] ),
    .B(_0416_),
    .X(_1330_));
 sky130_fd_sc_hd__xor2_1 _2595_ (.A(\transfer_count[2][22] ),
    .B(_0405_),
    .X(_1336_));
 sky130_fd_sc_hd__xnor2_1 _2596_ (.A(\transfer_count[2][20] ),
    .B(_0396_),
    .Y(_1342_));
 sky130_fd_sc_hd__xor2_1 _2597_ (.A(\transfer_count[2][18] ),
    .B(_0388_),
    .X(_1348_));
 sky130_fd_sc_hd__xor2_1 _2598_ (.A(\transfer_count[2][17] ),
    .B(_0383_),
    .X(_1351_));
 sky130_fd_sc_hd__xor2_1 _2599_ (.A(\transfer_count[2][16] ),
    .B(_0380_),
    .X(_1354_));
 sky130_fd_sc_hd__xor2_2 _2600_ (.A(\transfer_count[2][14] ),
    .B(_0366_),
    .X(_1360_));
 sky130_fd_sc_hd__xnor2_1 _2601_ (.A(\transfer_count[2][12] ),
    .B(_0357_),
    .Y(_1366_));
 sky130_fd_sc_hd__xor2_1 _2602_ (.A(_0347_),
    .B(_0349_),
    .X(_1372_));
 sky130_fd_sc_hd__xor2_2 _2603_ (.A(\transfer_count[2][8] ),
    .B(_0341_),
    .X(_1378_));
 sky130_fd_sc_hd__xnor2_1 _2604_ (.A(\transfer_count[2][6] ),
    .B(_0331_),
    .Y(_1384_));
 sky130_fd_sc_hd__xnor2_1 _2605_ (.A(\transfer_count[2][2] ),
    .B(_1399_),
    .Y(_1396_));
 sky130_fd_sc_hd__xor2_1 _2606_ (.A(\transfer_count[1][3] ),
    .B(_0460_),
    .X(_1417_));
 sky130_fd_sc_hd__xnor2_1 _2607_ (.A(_1412_),
    .B(\transfer_count[1][2] ),
    .Y(_1420_));
 sky130_fd_sc_hd__xor2_1 _2608_ (.A(\transfer_count[1][7] ),
    .B(_0473_),
    .X(_1423_));
 sky130_fd_sc_hd__xnor2_1 _2609_ (.A(_0800_),
    .B(_0468_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _2610_ (.A(_0553_),
    .B(_0554_),
    .Y(_0795_));
 sky130_fd_sc_hd__o21ai_1 _2611_ (.A1(_0553_),
    .A2(_0684_),
    .B1(_0795_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21o_1 _2612_ (.A1(_0445_),
    .A2(_0827_),
    .B1(_0695_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ai_0 _2613_ (.A1(_0671_),
    .A2(_0301_),
    .B1(_0701_),
    .Y(_0143_));
 sky130_fd_sc_hd__a21o_1 _2614_ (.A1(_0920_),
    .A2(_0921_),
    .B1(_0769_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2b_1 _2615_ (.A_N(net145),
    .B(_0666_),
    .Y(_0796_));
 sky130_fd_sc_hd__a21oi_1 _2616_ (.A1(_0667_),
    .A2(_0796_),
    .B1(_0920_),
    .Y(_0145_));
 sky130_fd_sc_hd__ha_1 _2617_ (.A(net75),
    .B(_1033_),
    .COUT(_1034_),
    .SUM(_1035_));
 sky130_fd_sc_hd__ha_1 _2618_ (.A(net74),
    .B(_1036_),
    .COUT(_1037_),
    .SUM(_1038_));
 sky130_fd_sc_hd__ha_1 _2619_ (.A(net73),
    .B(_1039_),
    .COUT(_1040_),
    .SUM(_1041_));
 sky130_fd_sc_hd__ha_1 _2620_ (.A(net72),
    .B(_1042_),
    .COUT(_1043_),
    .SUM(_1044_));
 sky130_fd_sc_hd__ha_1 _2621_ (.A(net71),
    .B(_1045_),
    .COUT(_1046_),
    .SUM(_1047_));
 sky130_fd_sc_hd__ha_1 _2622_ (.A(net70),
    .B(_1048_),
    .COUT(_1049_),
    .SUM(_1050_));
 sky130_fd_sc_hd__ha_1 _2623_ (.A(net69),
    .B(_1051_),
    .COUT(_1052_),
    .SUM(_1053_));
 sky130_fd_sc_hd__ha_1 _2624_ (.A(net68),
    .B(_1054_),
    .COUT(_1055_),
    .SUM(_1056_));
 sky130_fd_sc_hd__ha_1 _2625_ (.A(net93),
    .B(_1057_),
    .COUT(_1058_),
    .SUM(_1059_));
 sky130_fd_sc_hd__ha_1 _2626_ (.A(net92),
    .B(_1060_),
    .COUT(_1061_),
    .SUM(_1062_));
 sky130_fd_sc_hd__ha_1 _2627_ (.A(net91),
    .B(_1063_),
    .COUT(_1064_),
    .SUM(_1065_));
 sky130_fd_sc_hd__ha_1 _2628_ (.A(net90),
    .B(_1066_),
    .COUT(_1067_),
    .SUM(_1068_));
 sky130_fd_sc_hd__ha_1 _2629_ (.A(net88),
    .B(_1069_),
    .COUT(_1070_),
    .SUM(_1071_));
 sky130_fd_sc_hd__ha_1 _2630_ (.A(net87),
    .B(_1072_),
    .COUT(_1073_),
    .SUM(_1074_));
 sky130_fd_sc_hd__ha_1 _2631_ (.A(net86),
    .B(_1075_),
    .COUT(_1076_),
    .SUM(_1077_));
 sky130_fd_sc_hd__ha_1 _2632_ (.A(net85),
    .B(_1078_),
    .COUT(_1079_),
    .SUM(_1080_));
 sky130_fd_sc_hd__ha_1 _2633_ (.A(net84),
    .B(_1081_),
    .COUT(_1082_),
    .SUM(_1083_));
 sky130_fd_sc_hd__ha_1 _2634_ (.A(net83),
    .B(_1084_),
    .COUT(_1085_),
    .SUM(_1086_));
 sky130_fd_sc_hd__ha_1 _2635_ (.A(net82),
    .B(_1087_),
    .COUT(_1088_),
    .SUM(_1089_));
 sky130_fd_sc_hd__ha_1 _2636_ (.A(net81),
    .B(_1090_),
    .COUT(_1091_),
    .SUM(_1092_));
 sky130_fd_sc_hd__ha_1 _2637_ (.A(net80),
    .B(_1093_),
    .COUT(_1094_),
    .SUM(_1095_));
 sky130_fd_sc_hd__ha_1 _2638_ (.A(net79),
    .B(_1096_),
    .COUT(_1097_),
    .SUM(_1098_));
 sky130_fd_sc_hd__ha_1 _2639_ (.A(net77),
    .B(_1099_),
    .COUT(_1100_),
    .SUM(_1101_));
 sky130_fd_sc_hd__ha_1 _2640_ (.A(net76),
    .B(_1102_),
    .COUT(_1103_),
    .SUM(_1104_));
 sky130_fd_sc_hd__ha_1 _2641_ (.A(net36),
    .B(_1105_),
    .COUT(_1106_),
    .SUM(_1107_));
 sky130_fd_sc_hd__ha_1 _2642_ (.A(net35),
    .B(_1108_),
    .COUT(_1109_),
    .SUM(_1110_));
 sky130_fd_sc_hd__ha_1 _2643_ (.A(net34),
    .B(_1111_),
    .COUT(_1112_),
    .SUM(_1113_));
 sky130_fd_sc_hd__ha_1 _2644_ (.A(net33),
    .B(_1114_),
    .COUT(_1115_),
    .SUM(_1116_));
 sky130_fd_sc_hd__ha_1 _2645_ (.A(net32),
    .B(_1117_),
    .COUT(_1118_),
    .SUM(_1119_));
 sky130_fd_sc_hd__ha_1 _2646_ (.A(net31),
    .B(_1120_),
    .COUT(_1121_),
    .SUM(_1122_));
 sky130_fd_sc_hd__ha_1 _2647_ (.A(net30),
    .B(_1123_),
    .COUT(_1124_),
    .SUM(_1125_));
 sky130_fd_sc_hd__ha_1 _2648_ (.A(net29),
    .B(_1126_),
    .COUT(_1127_),
    .SUM(_1128_));
 sky130_fd_sc_hd__ha_1 _2649_ (.A(net27),
    .B(_1129_),
    .COUT(_1130_),
    .SUM(_1131_));
 sky130_fd_sc_hd__ha_1 _2650_ (.A(net26),
    .B(_1132_),
    .COUT(_1133_),
    .SUM(_1134_));
 sky130_fd_sc_hd__ha_1 _2651_ (.A(net25),
    .B(_1135_),
    .COUT(_1136_),
    .SUM(_1137_));
 sky130_fd_sc_hd__ha_1 _2652_ (.A(net24),
    .B(_1138_),
    .COUT(_1139_),
    .SUM(_1140_));
 sky130_fd_sc_hd__ha_1 _2653_ (.A(net23),
    .B(_1141_),
    .COUT(_1142_),
    .SUM(_1143_));
 sky130_fd_sc_hd__ha_1 _2654_ (.A(net22),
    .B(_1144_),
    .COUT(_1145_),
    .SUM(_1146_));
 sky130_fd_sc_hd__ha_1 _2655_ (.A(net21),
    .B(_1147_),
    .COUT(_1148_),
    .SUM(_1149_));
 sky130_fd_sc_hd__ha_1 _2656_ (.A(net20),
    .B(_1150_),
    .COUT(_1151_),
    .SUM(_1152_));
 sky130_fd_sc_hd__ha_1 _2657_ (.A(net19),
    .B(_1153_),
    .COUT(_1154_),
    .SUM(_1155_));
 sky130_fd_sc_hd__ha_1 _2658_ (.A(net18),
    .B(_1156_),
    .COUT(_1157_),
    .SUM(_1158_));
 sky130_fd_sc_hd__ha_1 _2659_ (.A(net16),
    .B(_1159_),
    .COUT(_1160_),
    .SUM(_1161_));
 sky130_fd_sc_hd__ha_1 _2660_ (.A(net15),
    .B(_1162_),
    .COUT(_1163_),
    .SUM(_1164_));
 sky130_fd_sc_hd__ha_1 _2661_ (.A(net14),
    .B(_1165_),
    .COUT(_1166_),
    .SUM(_1167_));
 sky130_fd_sc_hd__ha_1 _2662_ (.A(net13),
    .B(_1168_),
    .COUT(_1169_),
    .SUM(_1170_));
 sky130_fd_sc_hd__ha_1 _2663_ (.A(net12),
    .B(_1171_),
    .COUT(_1172_),
    .SUM(_1173_));
 sky130_fd_sc_hd__ha_1 _2664_ (.A(net11),
    .B(_1174_),
    .COUT(_1175_),
    .SUM(_1176_));
 sky130_fd_sc_hd__ha_1 _2665_ (.A(net10),
    .B(_1177_),
    .COUT(_1178_),
    .SUM(_1179_));
 sky130_fd_sc_hd__ha_1 _2666_ (.A(net9),
    .B(_1180_),
    .COUT(_1181_),
    .SUM(_1182_));
 sky130_fd_sc_hd__ha_1 _2667_ (.A(net8),
    .B(_1183_),
    .COUT(_1184_),
    .SUM(_1185_));
 sky130_fd_sc_hd__ha_1 _2668_ (.A(net7),
    .B(_1186_),
    .COUT(_1187_),
    .SUM(_1188_));
 sky130_fd_sc_hd__ha_1 _2669_ (.A(net132),
    .B(_1189_),
    .COUT(_1190_),
    .SUM(_1191_));
 sky130_fd_sc_hd__ha_1 _2670_ (.A(net131),
    .B(_1192_),
    .COUT(_1193_),
    .SUM(_1194_));
 sky130_fd_sc_hd__ha_1 _2671_ (.A(\transfer_count[3][0] ),
    .B(\transfer_count[3][1] ),
    .COUT(_1195_),
    .SUM(_1196_));
 sky130_fd_sc_hd__ha_1 _2672_ (.A(net130),
    .B(_1197_),
    .COUT(_1198_),
    .SUM(_1199_));
 sky130_fd_sc_hd__ha_1 _2673_ (.A(_1200_),
    .B(_1201_),
    .COUT(_1202_),
    .SUM(_1203_));
 sky130_fd_sc_hd__ha_1 _2674_ (.A(_1204_),
    .B(_1205_),
    .COUT(_1206_),
    .SUM(_1207_));
 sky130_fd_sc_hd__ha_2 _2675_ (.A(\transfer_count[0][0] ),
    .B(\transfer_count[0][1] ),
    .COUT(_1208_),
    .SUM(_1209_));
 sky130_fd_sc_hd__ha_1 _2676_ (.A(net45),
    .B(_1210_),
    .COUT(_1211_),
    .SUM(_1212_));
 sky130_fd_sc_hd__ha_1 _2677_ (.A(net67),
    .B(_1213_),
    .COUT(_1214_),
    .SUM(_1215_));
 sky130_fd_sc_hd__ha_1 _2678_ (.A(net56),
    .B(_1216_),
    .COUT(_1217_),
    .SUM(_1218_));
 sky130_fd_sc_hd__ha_1 _2679_ (.A(net111),
    .B(_1219_),
    .COUT(_1220_),
    .SUM(_1221_));
 sky130_fd_sc_hd__ha_1 _2680_ (.A(net100),
    .B(_1222_),
    .COUT(_1223_),
    .SUM(_1224_));
 sky130_fd_sc_hd__ha_1 _2681_ (.A(net89),
    .B(_1225_),
    .COUT(_1226_),
    .SUM(_1227_));
 sky130_fd_sc_hd__ha_1 _2682_ (.A(net78),
    .B(_1228_),
    .COUT(_1229_),
    .SUM(_1230_));
 sky130_fd_sc_hd__ha_1 _2683_ (.A(net40),
    .B(_1231_),
    .COUT(_1232_),
    .SUM(_1233_));
 sky130_fd_sc_hd__ha_1 _2684_ (.A(net39),
    .B(_1234_),
    .COUT(_1235_),
    .SUM(_1236_));
 sky130_fd_sc_hd__ha_1 _2685_ (.A(net38),
    .B(_1237_),
    .COUT(_1238_),
    .SUM(_1239_));
 sky130_fd_sc_hd__ha_1 _2686_ (.A(net37),
    .B(_1240_),
    .COUT(_1241_),
    .SUM(_1242_));
 sky130_fd_sc_hd__ha_1 _2687_ (.A(net28),
    .B(_1243_),
    .COUT(_1244_),
    .SUM(_1245_));
 sky130_fd_sc_hd__ha_1 _2688_ (.A(net17),
    .B(_1246_),
    .COUT(_1247_),
    .SUM(_1248_));
 sky130_fd_sc_hd__ha_1 _2689_ (.A(net133),
    .B(_1249_),
    .COUT(_1250_),
    .SUM(_1251_));
 sky130_fd_sc_hd__ha_1 _2690_ (.A(net122),
    .B(_1252_),
    .COUT(_1253_),
    .SUM(_1254_));
 sky130_fd_sc_hd__ha_1 _2691_ (.A(net58),
    .B(_1255_),
    .COUT(_1256_),
    .SUM(_1257_));
 sky130_fd_sc_hd__ha_1 _2692_ (.A(net57),
    .B(_1258_),
    .COUT(_1259_),
    .SUM(_1260_));
 sky130_fd_sc_hd__ha_1 _2693_ (.A(net55),
    .B(_1261_),
    .COUT(_1262_),
    .SUM(_1263_));
 sky130_fd_sc_hd__ha_1 _2694_ (.A(net54),
    .B(_1264_),
    .COUT(_1265_),
    .SUM(_1266_));
 sky130_fd_sc_hd__ha_1 _2695_ (.A(net53),
    .B(_1267_),
    .COUT(_1268_),
    .SUM(_1269_));
 sky130_fd_sc_hd__ha_1 _2696_ (.A(net52),
    .B(_1270_),
    .COUT(_1271_),
    .SUM(_1272_));
 sky130_fd_sc_hd__ha_1 _2697_ (.A(net51),
    .B(_1273_),
    .COUT(_1274_),
    .SUM(_1275_));
 sky130_fd_sc_hd__ha_1 _2698_ (.A(net50),
    .B(_1276_),
    .COUT(_1277_),
    .SUM(_1278_));
 sky130_fd_sc_hd__ha_1 _2699_ (.A(net49),
    .B(_1279_),
    .COUT(_1280_),
    .SUM(_1281_));
 sky130_fd_sc_hd__ha_1 _2700_ (.A(net48),
    .B(_1282_),
    .COUT(_1283_),
    .SUM(_1284_));
 sky130_fd_sc_hd__ha_1 _2701_ (.A(net47),
    .B(_1285_),
    .COUT(_1286_),
    .SUM(_1287_));
 sky130_fd_sc_hd__ha_1 _2702_ (.A(net46),
    .B(_1288_),
    .COUT(_1289_),
    .SUM(_1290_));
 sky130_fd_sc_hd__ha_1 _2703_ (.A(net44),
    .B(_1291_),
    .COUT(_1292_),
    .SUM(_1293_));
 sky130_fd_sc_hd__ha_1 _2704_ (.A(net43),
    .B(_1294_),
    .COUT(_1295_),
    .SUM(_1296_));
 sky130_fd_sc_hd__ha_1 _2705_ (.A(net42),
    .B(_1297_),
    .COUT(_1298_),
    .SUM(_1299_));
 sky130_fd_sc_hd__ha_1 _2706_ (.A(net41),
    .B(_1300_),
    .COUT(_1301_),
    .SUM(_1302_));
 sky130_fd_sc_hd__ha_1 _2707_ (.A(_1303_),
    .B(_1304_),
    .COUT(_1305_),
    .SUM(_1306_));
 sky130_fd_sc_hd__ha_1 _2708_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[1] ),
    .COUT(_1307_),
    .SUM(_1308_));
 sky130_fd_sc_hd__ha_1 _2709_ (.A(net128),
    .B(_1309_),
    .COUT(_1310_),
    .SUM(_1311_));
 sky130_fd_sc_hd__ha_1 _2710_ (.A(_1312_),
    .B(net127),
    .COUT(_1313_),
    .SUM(_1314_));
 sky130_fd_sc_hd__ha_1 _2711_ (.A(_1315_),
    .B(net126),
    .COUT(_1316_),
    .SUM(_1317_));
 sky130_fd_sc_hd__ha_1 _2712_ (.A(net125),
    .B(_1318_),
    .COUT(_1319_),
    .SUM(_1320_));
 sky130_fd_sc_hd__ha_1 _2713_ (.A(_1321_),
    .B(net124),
    .COUT(_1322_),
    .SUM(_1323_));
 sky130_fd_sc_hd__ha_1 _2714_ (.A(_1324_),
    .B(net123),
    .COUT(_1325_),
    .SUM(_1326_));
 sky130_fd_sc_hd__ha_1 _2715_ (.A(net121),
    .B(_1327_),
    .COUT(_1328_),
    .SUM(_1329_));
 sky130_fd_sc_hd__ha_1 _2716_ (.A(net120),
    .B(_1330_),
    .COUT(_1331_),
    .SUM(_1332_));
 sky130_fd_sc_hd__ha_1 _2717_ (.A(net119),
    .B(_1333_),
    .COUT(_1334_),
    .SUM(_1335_));
 sky130_fd_sc_hd__ha_1 _2718_ (.A(net118),
    .B(_1336_),
    .COUT(_1337_),
    .SUM(_1338_));
 sky130_fd_sc_hd__ha_1 _2719_ (.A(net117),
    .B(_1339_),
    .COUT(_1340_),
    .SUM(_1341_));
 sky130_fd_sc_hd__ha_1 _2720_ (.A(net116),
    .B(_1342_),
    .COUT(_1343_),
    .SUM(_1344_));
 sky130_fd_sc_hd__ha_1 _2721_ (.A(net115),
    .B(_1345_),
    .COUT(_1346_),
    .SUM(_1347_));
 sky130_fd_sc_hd__ha_1 _2722_ (.A(net114),
    .B(_1348_),
    .COUT(_1349_),
    .SUM(_1350_));
 sky130_fd_sc_hd__ha_1 _2723_ (.A(net113),
    .B(_1351_),
    .COUT(_1352_),
    .SUM(_1353_));
 sky130_fd_sc_hd__ha_1 _2724_ (.A(net112),
    .B(_1354_),
    .COUT(_1355_),
    .SUM(_1356_));
 sky130_fd_sc_hd__ha_1 _2725_ (.A(net110),
    .B(_1357_),
    .COUT(_1358_),
    .SUM(_1359_));
 sky130_fd_sc_hd__ha_1 _2726_ (.A(net109),
    .B(_1360_),
    .COUT(_1361_),
    .SUM(_1362_));
 sky130_fd_sc_hd__ha_1 _2727_ (.A(net108),
    .B(_1363_),
    .COUT(_1364_),
    .SUM(_1365_));
 sky130_fd_sc_hd__ha_1 _2728_ (.A(net107),
    .B(_1366_),
    .COUT(_1367_),
    .SUM(_1368_));
 sky130_fd_sc_hd__ha_1 _2729_ (.A(net106),
    .B(_1369_),
    .COUT(_1370_),
    .SUM(_1371_));
 sky130_fd_sc_hd__ha_1 _2730_ (.A(net105),
    .B(_1372_),
    .COUT(_1373_),
    .SUM(_1374_));
 sky130_fd_sc_hd__ha_1 _2731_ (.A(net104),
    .B(_1375_),
    .COUT(_1376_),
    .SUM(_1377_));
 sky130_fd_sc_hd__ha_1 _2732_ (.A(net103),
    .B(_1378_),
    .COUT(_1379_),
    .SUM(_1380_));
 sky130_fd_sc_hd__ha_1 _2733_ (.A(net102),
    .B(_1381_),
    .COUT(_1382_),
    .SUM(_1383_));
 sky130_fd_sc_hd__ha_1 _2734_ (.A(net101),
    .B(_1384_),
    .COUT(_1385_),
    .SUM(_1386_));
 sky130_fd_sc_hd__ha_1 _2735_ (.A(net99),
    .B(_1387_),
    .COUT(_1388_),
    .SUM(_1389_));
 sky130_fd_sc_hd__ha_1 _2736_ (.A(net98),
    .B(_1390_),
    .COUT(_1391_),
    .SUM(_1392_));
 sky130_fd_sc_hd__ha_1 _2737_ (.A(net97),
    .B(_1393_),
    .COUT(_1394_),
    .SUM(_1395_));
 sky130_fd_sc_hd__ha_1 _2738_ (.A(net96),
    .B(_1396_),
    .COUT(_1397_),
    .SUM(_1398_));
 sky130_fd_sc_hd__ha_1 _2739_ (.A(\transfer_count[2][0] ),
    .B(\transfer_count[2][1] ),
    .COUT(_1399_),
    .SUM(_1400_));
 sky130_fd_sc_hd__ha_1 _2740_ (.A(net95),
    .B(_1401_),
    .COUT(_1402_),
    .SUM(_1403_));
 sky130_fd_sc_hd__ha_1 _2741_ (.A(_1404_),
    .B(_1405_),
    .COUT(_1406_),
    .SUM(_1407_));
 sky130_fd_sc_hd__ha_1 _2742_ (.A(_1408_),
    .B(_1409_),
    .COUT(_1410_),
    .SUM(_1411_));
 sky130_fd_sc_hd__ha_1 _2743_ (.A(\transfer_count[1][0] ),
    .B(\transfer_count[1][1] ),
    .COUT(_1412_),
    .SUM(_1413_));
 sky130_fd_sc_hd__ha_1 _2744_ (.A(net60),
    .B(_1414_),
    .COUT(_1415_),
    .SUM(_1416_));
 sky130_fd_sc_hd__ha_1 _2745_ (.A(net62),
    .B(_1417_),
    .COUT(_1418_),
    .SUM(_1419_));
 sky130_fd_sc_hd__ha_1 _2746_ (.A(net61),
    .B(_1420_),
    .COUT(_1421_),
    .SUM(_1422_));
 sky130_fd_sc_hd__ha_1 _2747_ (.A(net66),
    .B(_1423_),
    .COUT(_1424_),
    .SUM(_1425_));
 sky130_fd_sc_hd__ha_1 _2748_ (.A(net65),
    .B(_1426_),
    .COUT(_1427_),
    .SUM(_1428_));
 sky130_fd_sc_hd__ha_1 _2749_ (.A(net64),
    .B(_1429_),
    .COUT(_1430_),
    .SUM(_1431_));
 sky130_fd_sc_hd__ha_1 _2750_ (.A(net63),
    .B(_1432_),
    .COUT(_1433_),
    .SUM(_1434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 _2752_ (.A(net175),
    .X(debug_channel_state[0]));
 sky130_fd_sc_hd__buf_4 _2753_ (.A(net176),
    .X(debug_channel_state[1]));
 sky130_fd_sc_hd__buf_4 _2754_ (.A(net177),
    .X(debug_channel_state[2]));
 sky130_fd_sc_hd__buf_4 _2755_ (.A(net178),
    .X(debug_channel_state[3]));
 sky130_fd_sc_hd__buf_4 _2756_ (.A(net179),
    .X(debug_channel_state[4]));
 sky130_fd_sc_hd__buf_4 _2757_ (.A(net180),
    .X(debug_channel_state[5]));
 sky130_fd_sc_hd__buf_4 _2758_ (.A(net181),
    .X(debug_channel_state[6]));
 sky130_fd_sc_hd__buf_4 _2759_ (.A(net182),
    .X(debug_channel_state[7]));
 sky130_fd_sc_hd__buf_4 _2760_ (.A(net183),
    .X(debug_channel_state[8]));
 sky130_fd_sc_hd__buf_4 _2761_ (.A(net184),
    .X(debug_channel_state[9]));
 sky130_fd_sc_hd__buf_4 _2762_ (.A(net185),
    .X(debug_channel_state[10]));
 sky130_fd_sc_hd__buf_4 _2763_ (.A(net186),
    .X(debug_channel_state[11]));
 sky130_fd_sc_hd__buf_4 _2764_ (.A(net187),
    .X(debug_transfer_count[0]));
 sky130_fd_sc_hd__buf_4 _2765_ (.A(net188),
    .X(debug_transfer_count[1]));
 sky130_fd_sc_hd__buf_4 _2766_ (.A(net189),
    .X(debug_transfer_count[2]));
 sky130_fd_sc_hd__buf_4 _2767_ (.A(net190),
    .X(debug_transfer_count[3]));
 sky130_fd_sc_hd__buf_4 _2768_ (.A(net191),
    .X(debug_transfer_count[4]));
 sky130_fd_sc_hd__buf_4 _2769_ (.A(net192),
    .X(debug_transfer_count[5]));
 sky130_fd_sc_hd__buf_4 _2770_ (.A(net193),
    .X(debug_transfer_count[6]));
 sky130_fd_sc_hd__buf_4 _2771_ (.A(net194),
    .X(debug_transfer_count[7]));
 sky130_fd_sc_hd__buf_4 _2772_ (.A(net195),
    .X(debug_transfer_count[8]));
 sky130_fd_sc_hd__buf_4 _2773_ (.A(net196),
    .X(debug_transfer_count[9]));
 sky130_fd_sc_hd__buf_4 _2774_ (.A(net197),
    .X(debug_transfer_count[10]));
 sky130_fd_sc_hd__buf_4 _2775_ (.A(net198),
    .X(debug_transfer_count[11]));
 sky130_fd_sc_hd__buf_4 _2776_ (.A(net199),
    .X(debug_transfer_count[12]));
 sky130_fd_sc_hd__buf_4 _2777_ (.A(net200),
    .X(debug_transfer_count[13]));
 sky130_fd_sc_hd__buf_4 _2778_ (.A(net201),
    .X(debug_transfer_count[14]));
 sky130_fd_sc_hd__buf_4 _2779_ (.A(net202),
    .X(debug_transfer_count[15]));
 sky130_fd_sc_hd__buf_4 _2780_ (.A(net203),
    .X(debug_transfer_count[16]));
 sky130_fd_sc_hd__buf_4 _2781_ (.A(net204),
    .X(debug_transfer_count[17]));
 sky130_fd_sc_hd__buf_4 _2782_ (.A(net205),
    .X(debug_transfer_count[18]));
 sky130_fd_sc_hd__buf_4 _2783_ (.A(net206),
    .X(debug_transfer_count[19]));
 sky130_fd_sc_hd__buf_4 _2784_ (.A(net207),
    .X(debug_transfer_count[20]));
 sky130_fd_sc_hd__buf_4 _2785_ (.A(net208),
    .X(debug_transfer_count[21]));
 sky130_fd_sc_hd__buf_4 _2786_ (.A(net209),
    .X(debug_transfer_count[22]));
 sky130_fd_sc_hd__buf_4 _2787_ (.A(net210),
    .X(debug_transfer_count[23]));
 sky130_fd_sc_hd__buf_4 _2788_ (.A(net211),
    .X(debug_transfer_count[24]));
 sky130_fd_sc_hd__buf_4 _2789_ (.A(net212),
    .X(debug_transfer_count[25]));
 sky130_fd_sc_hd__buf_4 _2790_ (.A(net213),
    .X(debug_transfer_count[26]));
 sky130_fd_sc_hd__buf_4 _2791_ (.A(net214),
    .X(debug_transfer_count[27]));
 sky130_fd_sc_hd__buf_4 _2792_ (.A(net215),
    .X(debug_transfer_count[28]));
 sky130_fd_sc_hd__buf_4 _2793_ (.A(net216),
    .X(debug_transfer_count[29]));
 sky130_fd_sc_hd__buf_4 _2794_ (.A(net217),
    .X(debug_transfer_count[30]));
 sky130_fd_sc_hd__buf_4 _2795_ (.A(net218),
    .X(debug_transfer_count[31]));
 sky130_fd_sc_hd__buf_4 _2796_ (.A(net219),
    .X(debug_transfer_count[32]));
 sky130_fd_sc_hd__buf_4 _2797_ (.A(net220),
    .X(debug_transfer_count[33]));
 sky130_fd_sc_hd__buf_4 _2798_ (.A(net221),
    .X(debug_transfer_count[34]));
 sky130_fd_sc_hd__buf_4 _2799_ (.A(net222),
    .X(debug_transfer_count[35]));
 sky130_fd_sc_hd__buf_4 _2800_ (.A(net223),
    .X(debug_transfer_count[36]));
 sky130_fd_sc_hd__buf_4 _2801_ (.A(net224),
    .X(debug_transfer_count[37]));
 sky130_fd_sc_hd__buf_4 _2802_ (.A(net225),
    .X(debug_transfer_count[38]));
 sky130_fd_sc_hd__buf_4 _2803_ (.A(net226),
    .X(debug_transfer_count[39]));
 sky130_fd_sc_hd__buf_4 _2804_ (.A(net227),
    .X(debug_transfer_count[40]));
 sky130_fd_sc_hd__buf_4 _2805_ (.A(net228),
    .X(debug_transfer_count[41]));
 sky130_fd_sc_hd__buf_4 _2806_ (.A(net229),
    .X(debug_transfer_count[42]));
 sky130_fd_sc_hd__buf_4 _2807_ (.A(net230),
    .X(debug_transfer_count[43]));
 sky130_fd_sc_hd__buf_4 _2808_ (.A(net231),
    .X(debug_transfer_count[44]));
 sky130_fd_sc_hd__buf_4 _2809_ (.A(net232),
    .X(debug_transfer_count[45]));
 sky130_fd_sc_hd__buf_4 _2810_ (.A(net233),
    .X(debug_transfer_count[46]));
 sky130_fd_sc_hd__buf_4 _2811_ (.A(net234),
    .X(debug_transfer_count[47]));
 sky130_fd_sc_hd__buf_4 _2812_ (.A(net235),
    .X(debug_transfer_count[48]));
 sky130_fd_sc_hd__buf_4 _2813_ (.A(net236),
    .X(debug_transfer_count[49]));
 sky130_fd_sc_hd__buf_4 _2814_ (.A(net237),
    .X(debug_transfer_count[50]));
 sky130_fd_sc_hd__buf_4 _2815_ (.A(net238),
    .X(debug_transfer_count[51]));
 sky130_fd_sc_hd__buf_4 _2816_ (.A(net239),
    .X(debug_transfer_count[52]));
 sky130_fd_sc_hd__buf_4 _2817_ (.A(net240),
    .X(debug_transfer_count[53]));
 sky130_fd_sc_hd__buf_4 _2818_ (.A(net241),
    .X(debug_transfer_count[54]));
 sky130_fd_sc_hd__buf_4 _2819_ (.A(net242),
    .X(debug_transfer_count[55]));
 sky130_fd_sc_hd__buf_4 _2820_ (.A(net243),
    .X(debug_transfer_count[56]));
 sky130_fd_sc_hd__buf_4 _2821_ (.A(net244),
    .X(debug_transfer_count[57]));
 sky130_fd_sc_hd__buf_4 _2822_ (.A(net245),
    .X(debug_transfer_count[58]));
 sky130_fd_sc_hd__buf_4 _2823_ (.A(net246),
    .X(debug_transfer_count[59]));
 sky130_fd_sc_hd__buf_4 _2824_ (.A(net247),
    .X(debug_transfer_count[60]));
 sky130_fd_sc_hd__buf_4 _2825_ (.A(net248),
    .X(debug_transfer_count[61]));
 sky130_fd_sc_hd__buf_4 _2826_ (.A(net249),
    .X(debug_transfer_count[62]));
 sky130_fd_sc_hd__buf_4 _2827_ (.A(net250),
    .X(debug_transfer_count[63]));
 sky130_fd_sc_hd__buf_4 _2828_ (.A(net251),
    .X(debug_transfer_count[64]));
 sky130_fd_sc_hd__buf_4 _2829_ (.A(net252),
    .X(debug_transfer_count[65]));
 sky130_fd_sc_hd__buf_4 _2830_ (.A(net253),
    .X(debug_transfer_count[66]));
 sky130_fd_sc_hd__buf_4 _2831_ (.A(net254),
    .X(debug_transfer_count[67]));
 sky130_fd_sc_hd__buf_4 _2832_ (.A(net255),
    .X(debug_transfer_count[68]));
 sky130_fd_sc_hd__buf_4 _2833_ (.A(net256),
    .X(debug_transfer_count[69]));
 sky130_fd_sc_hd__buf_4 _2834_ (.A(net257),
    .X(debug_transfer_count[70]));
 sky130_fd_sc_hd__buf_4 _2835_ (.A(net258),
    .X(debug_transfer_count[71]));
 sky130_fd_sc_hd__buf_4 _2836_ (.A(net259),
    .X(debug_transfer_count[72]));
 sky130_fd_sc_hd__buf_4 _2837_ (.A(net260),
    .X(debug_transfer_count[73]));
 sky130_fd_sc_hd__buf_4 _2838_ (.A(net261),
    .X(debug_transfer_count[74]));
 sky130_fd_sc_hd__buf_4 _2839_ (.A(net262),
    .X(debug_transfer_count[75]));
 sky130_fd_sc_hd__buf_4 _2840_ (.A(net263),
    .X(debug_transfer_count[76]));
 sky130_fd_sc_hd__buf_4 _2841_ (.A(net264),
    .X(debug_transfer_count[77]));
 sky130_fd_sc_hd__buf_4 _2842_ (.A(net265),
    .X(debug_transfer_count[78]));
 sky130_fd_sc_hd__buf_4 _2843_ (.A(net266),
    .X(debug_transfer_count[79]));
 sky130_fd_sc_hd__buf_4 _2844_ (.A(net267),
    .X(debug_transfer_count[80]));
 sky130_fd_sc_hd__buf_4 _2845_ (.A(net268),
    .X(debug_transfer_count[81]));
 sky130_fd_sc_hd__buf_4 _2846_ (.A(net269),
    .X(debug_transfer_count[82]));
 sky130_fd_sc_hd__buf_4 _2847_ (.A(net270),
    .X(debug_transfer_count[83]));
 sky130_fd_sc_hd__buf_4 _2848_ (.A(net271),
    .X(debug_transfer_count[84]));
 sky130_fd_sc_hd__buf_4 _2849_ (.A(net272),
    .X(debug_transfer_count[85]));
 sky130_fd_sc_hd__buf_4 _2850_ (.A(net273),
    .X(debug_transfer_count[86]));
 sky130_fd_sc_hd__buf_4 _2851_ (.A(net274),
    .X(debug_transfer_count[87]));
 sky130_fd_sc_hd__buf_4 _2852_ (.A(net275),
    .X(debug_transfer_count[88]));
 sky130_fd_sc_hd__buf_4 _2853_ (.A(net276),
    .X(debug_transfer_count[89]));
 sky130_fd_sc_hd__buf_4 _2854_ (.A(net277),
    .X(debug_transfer_count[90]));
 sky130_fd_sc_hd__buf_4 _2855_ (.A(net278),
    .X(debug_transfer_count[91]));
 sky130_fd_sc_hd__buf_4 _2856_ (.A(net279),
    .X(debug_transfer_count[92]));
 sky130_fd_sc_hd__buf_4 _2857_ (.A(net280),
    .X(debug_transfer_count[93]));
 sky130_fd_sc_hd__buf_4 _2858_ (.A(net281),
    .X(debug_transfer_count[94]));
 sky130_fd_sc_hd__buf_4 _2859_ (.A(net282),
    .X(debug_transfer_count[95]));
 sky130_fd_sc_hd__buf_4 _2860_ (.A(net283),
    .X(debug_transfer_count[96]));
 sky130_fd_sc_hd__buf_4 _2861_ (.A(net284),
    .X(debug_transfer_count[97]));
 sky130_fd_sc_hd__buf_4 _2862_ (.A(net285),
    .X(debug_transfer_count[98]));
 sky130_fd_sc_hd__buf_4 _2863_ (.A(net286),
    .X(debug_transfer_count[99]));
 sky130_fd_sc_hd__buf_4 _2864_ (.A(net287),
    .X(debug_transfer_count[100]));
 sky130_fd_sc_hd__buf_4 _2865_ (.A(net288),
    .X(debug_transfer_count[101]));
 sky130_fd_sc_hd__buf_4 _2866_ (.A(net289),
    .X(debug_transfer_count[102]));
 sky130_fd_sc_hd__buf_4 _2867_ (.A(net290),
    .X(debug_transfer_count[103]));
 sky130_fd_sc_hd__buf_4 _2868_ (.A(net291),
    .X(debug_transfer_count[104]));
 sky130_fd_sc_hd__buf_4 _2869_ (.A(net292),
    .X(debug_transfer_count[105]));
 sky130_fd_sc_hd__buf_4 _2870_ (.A(net293),
    .X(debug_transfer_count[106]));
 sky130_fd_sc_hd__buf_4 _2871_ (.A(net294),
    .X(debug_transfer_count[107]));
 sky130_fd_sc_hd__buf_4 _2872_ (.A(net295),
    .X(debug_transfer_count[108]));
 sky130_fd_sc_hd__buf_4 _2873_ (.A(net296),
    .X(debug_transfer_count[109]));
 sky130_fd_sc_hd__buf_4 _2874_ (.A(net297),
    .X(debug_transfer_count[110]));
 sky130_fd_sc_hd__buf_4 _2875_ (.A(net298),
    .X(debug_transfer_count[111]));
 sky130_fd_sc_hd__buf_4 _2876_ (.A(net299),
    .X(debug_transfer_count[112]));
 sky130_fd_sc_hd__buf_4 _2877_ (.A(net300),
    .X(debug_transfer_count[113]));
 sky130_fd_sc_hd__buf_4 _2878_ (.A(net301),
    .X(debug_transfer_count[114]));
 sky130_fd_sc_hd__buf_4 _2879_ (.A(net302),
    .X(debug_transfer_count[115]));
 sky130_fd_sc_hd__buf_4 _2880_ (.A(net303),
    .X(debug_transfer_count[116]));
 sky130_fd_sc_hd__buf_4 _2881_ (.A(net304),
    .X(debug_transfer_count[117]));
 sky130_fd_sc_hd__buf_4 _2882_ (.A(net305),
    .X(debug_transfer_count[118]));
 sky130_fd_sc_hd__buf_4 _2883_ (.A(net306),
    .X(debug_transfer_count[119]));
 sky130_fd_sc_hd__buf_4 _2884_ (.A(net307),
    .X(debug_transfer_count[120]));
 sky130_fd_sc_hd__buf_4 _2885_ (.A(net308),
    .X(debug_transfer_count[121]));
 sky130_fd_sc_hd__buf_4 _2886_ (.A(net309),
    .X(debug_transfer_count[122]));
 sky130_fd_sc_hd__buf_4 _2887_ (.A(net310),
    .X(debug_transfer_count[123]));
 sky130_fd_sc_hd__buf_4 _2888_ (.A(net311),
    .X(debug_transfer_count[124]));
 sky130_fd_sc_hd__buf_4 _2889_ (.A(net312),
    .X(debug_transfer_count[125]));
 sky130_fd_sc_hd__buf_4 _2890_ (.A(net313),
    .X(debug_transfer_count[126]));
 sky130_fd_sc_hd__buf_4 _2891_ (.A(net314),
    .X(debug_transfer_count[127]));
 sky130_fd_sc_hd__buf_4 _2892_ (.A(net315),
    .X(dst_addr[0]));
 sky130_fd_sc_hd__buf_4 _2893_ (.A(net316),
    .X(dst_addr[1]));
 sky130_fd_sc_hd__buf_4 _2894_ (.A(net317),
    .X(dst_addr[2]));
 sky130_fd_sc_hd__buf_4 _2895_ (.A(net318),
    .X(dst_addr[3]));
 sky130_fd_sc_hd__buf_4 _2896_ (.A(net319),
    .X(dst_addr[4]));
 sky130_fd_sc_hd__buf_4 _2897_ (.A(net320),
    .X(dst_addr[5]));
 sky130_fd_sc_hd__buf_4 _2898_ (.A(net321),
    .X(dst_addr[6]));
 sky130_fd_sc_hd__buf_4 _2899_ (.A(net322),
    .X(dst_addr[7]));
 sky130_fd_sc_hd__buf_4 _2900_ (.A(net323),
    .X(dst_addr[8]));
 sky130_fd_sc_hd__buf_4 _2901_ (.A(net324),
    .X(dst_addr[9]));
 sky130_fd_sc_hd__buf_4 _2902_ (.A(net325),
    .X(dst_addr[10]));
 sky130_fd_sc_hd__buf_4 _2903_ (.A(net326),
    .X(dst_addr[11]));
 sky130_fd_sc_hd__buf_4 _2904_ (.A(net327),
    .X(dst_addr[12]));
 sky130_fd_sc_hd__buf_4 _2905_ (.A(net328),
    .X(dst_addr[13]));
 sky130_fd_sc_hd__buf_4 _2906_ (.A(net329),
    .X(dst_addr[14]));
 sky130_fd_sc_hd__buf_4 _2907_ (.A(net330),
    .X(dst_addr[15]));
 sky130_fd_sc_hd__buf_4 _2908_ (.A(net331),
    .X(dst_addr[16]));
 sky130_fd_sc_hd__buf_4 _2909_ (.A(net332),
    .X(dst_addr[17]));
 sky130_fd_sc_hd__buf_4 _2910_ (.A(net333),
    .X(dst_addr[18]));
 sky130_fd_sc_hd__buf_4 _2911_ (.A(net334),
    .X(dst_addr[19]));
 sky130_fd_sc_hd__buf_4 _2912_ (.A(net335),
    .X(dst_addr[20]));
 sky130_fd_sc_hd__buf_4 _2913_ (.A(net336),
    .X(dst_addr[21]));
 sky130_fd_sc_hd__buf_4 _2914_ (.A(net337),
    .X(dst_addr[22]));
 sky130_fd_sc_hd__buf_4 _2915_ (.A(net338),
    .X(dst_addr[23]));
 sky130_fd_sc_hd__buf_4 _2916_ (.A(net339),
    .X(dst_addr[24]));
 sky130_fd_sc_hd__buf_4 _2917_ (.A(net340),
    .X(dst_addr[25]));
 sky130_fd_sc_hd__buf_4 _2918_ (.A(net341),
    .X(dst_addr[26]));
 sky130_fd_sc_hd__buf_4 _2919_ (.A(net342),
    .X(dst_addr[27]));
 sky130_fd_sc_hd__buf_4 _2920_ (.A(net343),
    .X(dst_addr[28]));
 sky130_fd_sc_hd__buf_4 _2921_ (.A(net344),
    .X(dst_addr[29]));
 sky130_fd_sc_hd__buf_4 _2922_ (.A(net345),
    .X(dst_addr[30]));
 sky130_fd_sc_hd__buf_4 _2923_ (.A(net346),
    .X(dst_addr[31]));
 sky130_fd_sc_hd__buf_4 _2924_ (.A(net347),
    .X(dst_addr[32]));
 sky130_fd_sc_hd__buf_4 _2925_ (.A(net348),
    .X(dst_addr[33]));
 sky130_fd_sc_hd__buf_4 _2926_ (.A(net349),
    .X(dst_addr[34]));
 sky130_fd_sc_hd__buf_4 _2927_ (.A(net350),
    .X(dst_addr[35]));
 sky130_fd_sc_hd__buf_4 _2928_ (.A(net351),
    .X(dst_addr[36]));
 sky130_fd_sc_hd__buf_4 _2929_ (.A(net352),
    .X(dst_addr[37]));
 sky130_fd_sc_hd__buf_4 _2930_ (.A(net353),
    .X(dst_addr[38]));
 sky130_fd_sc_hd__buf_4 _2931_ (.A(net354),
    .X(dst_addr[39]));
 sky130_fd_sc_hd__buf_4 _2932_ (.A(net355),
    .X(dst_addr[40]));
 sky130_fd_sc_hd__buf_4 _2933_ (.A(net356),
    .X(dst_addr[41]));
 sky130_fd_sc_hd__buf_4 _2934_ (.A(net357),
    .X(dst_addr[42]));
 sky130_fd_sc_hd__buf_4 _2935_ (.A(net358),
    .X(dst_addr[43]));
 sky130_fd_sc_hd__buf_4 _2936_ (.A(net359),
    .X(dst_addr[44]));
 sky130_fd_sc_hd__buf_4 _2937_ (.A(net360),
    .X(dst_addr[45]));
 sky130_fd_sc_hd__buf_4 _2938_ (.A(net361),
    .X(dst_addr[46]));
 sky130_fd_sc_hd__buf_4 _2939_ (.A(net362),
    .X(dst_addr[47]));
 sky130_fd_sc_hd__buf_4 _2940_ (.A(net363),
    .X(dst_addr[48]));
 sky130_fd_sc_hd__buf_4 _2941_ (.A(net364),
    .X(dst_addr[49]));
 sky130_fd_sc_hd__buf_4 _2942_ (.A(net365),
    .X(dst_addr[50]));
 sky130_fd_sc_hd__buf_4 _2943_ (.A(net366),
    .X(dst_addr[51]));
 sky130_fd_sc_hd__buf_4 _2944_ (.A(net367),
    .X(dst_addr[52]));
 sky130_fd_sc_hd__buf_4 _2945_ (.A(net368),
    .X(dst_addr[53]));
 sky130_fd_sc_hd__buf_4 _2946_ (.A(net369),
    .X(dst_addr[54]));
 sky130_fd_sc_hd__buf_4 _2947_ (.A(net370),
    .X(dst_addr[55]));
 sky130_fd_sc_hd__buf_4 _2948_ (.A(net371),
    .X(dst_addr[56]));
 sky130_fd_sc_hd__buf_4 _2949_ (.A(net372),
    .X(dst_addr[57]));
 sky130_fd_sc_hd__buf_4 _2950_ (.A(net373),
    .X(dst_addr[58]));
 sky130_fd_sc_hd__buf_4 _2951_ (.A(net374),
    .X(dst_addr[59]));
 sky130_fd_sc_hd__buf_4 _2952_ (.A(net375),
    .X(dst_addr[60]));
 sky130_fd_sc_hd__buf_4 _2953_ (.A(net376),
    .X(dst_addr[61]));
 sky130_fd_sc_hd__buf_4 _2954_ (.A(net377),
    .X(dst_addr[62]));
 sky130_fd_sc_hd__buf_4 _2955_ (.A(net378),
    .X(dst_addr[63]));
 sky130_fd_sc_hd__buf_4 _2956_ (.A(net379),
    .X(dst_addr[64]));
 sky130_fd_sc_hd__buf_4 _2957_ (.A(net380),
    .X(dst_addr[65]));
 sky130_fd_sc_hd__buf_4 _2958_ (.A(net381),
    .X(dst_addr[66]));
 sky130_fd_sc_hd__buf_4 _2959_ (.A(net382),
    .X(dst_addr[67]));
 sky130_fd_sc_hd__buf_4 _2960_ (.A(net383),
    .X(dst_addr[68]));
 sky130_fd_sc_hd__buf_4 _2961_ (.A(net384),
    .X(dst_addr[69]));
 sky130_fd_sc_hd__buf_4 _2962_ (.A(net385),
    .X(dst_addr[70]));
 sky130_fd_sc_hd__buf_4 _2963_ (.A(net386),
    .X(dst_addr[71]));
 sky130_fd_sc_hd__buf_4 _2964_ (.A(net387),
    .X(dst_addr[72]));
 sky130_fd_sc_hd__buf_4 _2965_ (.A(net388),
    .X(dst_addr[73]));
 sky130_fd_sc_hd__buf_4 _2966_ (.A(net389),
    .X(dst_addr[74]));
 sky130_fd_sc_hd__buf_4 _2967_ (.A(net390),
    .X(dst_addr[75]));
 sky130_fd_sc_hd__buf_4 _2968_ (.A(net391),
    .X(dst_addr[76]));
 sky130_fd_sc_hd__buf_4 _2969_ (.A(net392),
    .X(dst_addr[77]));
 sky130_fd_sc_hd__buf_4 _2970_ (.A(net393),
    .X(dst_addr[78]));
 sky130_fd_sc_hd__buf_4 _2971_ (.A(net394),
    .X(dst_addr[79]));
 sky130_fd_sc_hd__buf_4 _2972_ (.A(net395),
    .X(dst_addr[80]));
 sky130_fd_sc_hd__buf_4 _2973_ (.A(net396),
    .X(dst_addr[81]));
 sky130_fd_sc_hd__buf_4 _2974_ (.A(net397),
    .X(dst_addr[82]));
 sky130_fd_sc_hd__buf_4 _2975_ (.A(net398),
    .X(dst_addr[83]));
 sky130_fd_sc_hd__buf_4 _2976_ (.A(net399),
    .X(dst_addr[84]));
 sky130_fd_sc_hd__buf_4 _2977_ (.A(net400),
    .X(dst_addr[85]));
 sky130_fd_sc_hd__buf_4 _2978_ (.A(net401),
    .X(dst_addr[86]));
 sky130_fd_sc_hd__buf_4 _2979_ (.A(net402),
    .X(dst_addr[87]));
 sky130_fd_sc_hd__buf_4 _2980_ (.A(net403),
    .X(dst_addr[88]));
 sky130_fd_sc_hd__buf_4 _2981_ (.A(net404),
    .X(dst_addr[89]));
 sky130_fd_sc_hd__buf_4 _2982_ (.A(net405),
    .X(dst_addr[90]));
 sky130_fd_sc_hd__buf_4 _2983_ (.A(net406),
    .X(dst_addr[91]));
 sky130_fd_sc_hd__buf_4 _2984_ (.A(net407),
    .X(dst_addr[92]));
 sky130_fd_sc_hd__buf_4 _2985_ (.A(net408),
    .X(dst_addr[93]));
 sky130_fd_sc_hd__buf_4 _2986_ (.A(net409),
    .X(dst_addr[94]));
 sky130_fd_sc_hd__buf_4 _2987_ (.A(net410),
    .X(dst_addr[95]));
 sky130_fd_sc_hd__buf_4 _2988_ (.A(net411),
    .X(dst_addr[96]));
 sky130_fd_sc_hd__buf_4 _2989_ (.A(net412),
    .X(dst_addr[97]));
 sky130_fd_sc_hd__buf_4 _2990_ (.A(net413),
    .X(dst_addr[98]));
 sky130_fd_sc_hd__buf_4 _2991_ (.A(net414),
    .X(dst_addr[99]));
 sky130_fd_sc_hd__buf_4 _2992_ (.A(net415),
    .X(dst_addr[100]));
 sky130_fd_sc_hd__buf_4 _2993_ (.A(net416),
    .X(dst_addr[101]));
 sky130_fd_sc_hd__buf_4 _2994_ (.A(net417),
    .X(dst_addr[102]));
 sky130_fd_sc_hd__buf_4 _2995_ (.A(net418),
    .X(dst_addr[103]));
 sky130_fd_sc_hd__buf_4 _2996_ (.A(net419),
    .X(dst_addr[104]));
 sky130_fd_sc_hd__buf_4 _2997_ (.A(net420),
    .X(dst_addr[105]));
 sky130_fd_sc_hd__buf_4 _2998_ (.A(net421),
    .X(dst_addr[106]));
 sky130_fd_sc_hd__buf_4 _2999_ (.A(net422),
    .X(dst_addr[107]));
 sky130_fd_sc_hd__buf_4 _3000_ (.A(net423),
    .X(dst_addr[108]));
 sky130_fd_sc_hd__buf_4 _3001_ (.A(net424),
    .X(dst_addr[109]));
 sky130_fd_sc_hd__buf_4 _3002_ (.A(net425),
    .X(dst_addr[110]));
 sky130_fd_sc_hd__buf_4 _3003_ (.A(net426),
    .X(dst_addr[111]));
 sky130_fd_sc_hd__buf_4 _3004_ (.A(net427),
    .X(dst_addr[112]));
 sky130_fd_sc_hd__buf_4 _3005_ (.A(net428),
    .X(dst_addr[113]));
 sky130_fd_sc_hd__buf_4 _3006_ (.A(net429),
    .X(dst_addr[114]));
 sky130_fd_sc_hd__buf_4 _3007_ (.A(net430),
    .X(dst_addr[115]));
 sky130_fd_sc_hd__buf_4 _3008_ (.A(net431),
    .X(dst_addr[116]));
 sky130_fd_sc_hd__buf_4 _3009_ (.A(net432),
    .X(dst_addr[117]));
 sky130_fd_sc_hd__buf_4 _3010_ (.A(net433),
    .X(dst_addr[118]));
 sky130_fd_sc_hd__buf_4 _3011_ (.A(net434),
    .X(dst_addr[119]));
 sky130_fd_sc_hd__buf_4 _3012_ (.A(net435),
    .X(dst_addr[120]));
 sky130_fd_sc_hd__buf_4 _3013_ (.A(net436),
    .X(dst_addr[121]));
 sky130_fd_sc_hd__buf_4 _3014_ (.A(net437),
    .X(dst_addr[122]));
 sky130_fd_sc_hd__buf_4 _3015_ (.A(net438),
    .X(dst_addr[123]));
 sky130_fd_sc_hd__buf_4 _3016_ (.A(net439),
    .X(dst_addr[124]));
 sky130_fd_sc_hd__buf_4 _3017_ (.A(net440),
    .X(dst_addr[125]));
 sky130_fd_sc_hd__buf_4 _3018_ (.A(net441),
    .X(dst_addr[126]));
 sky130_fd_sc_hd__buf_4 _3019_ (.A(net442),
    .X(dst_addr[127]));
 sky130_fd_sc_hd__buf_4 _3020_ (.A(net443),
    .X(dst_wdata[0]));
 sky130_fd_sc_hd__buf_4 _3021_ (.A(net444),
    .X(dst_wdata[1]));
 sky130_fd_sc_hd__buf_4 _3022_ (.A(net445),
    .X(dst_wdata[2]));
 sky130_fd_sc_hd__buf_4 _3023_ (.A(net446),
    .X(dst_wdata[3]));
 sky130_fd_sc_hd__buf_4 _3024_ (.A(net447),
    .X(dst_wdata[4]));
 sky130_fd_sc_hd__buf_4 _3025_ (.A(net448),
    .X(dst_wdata[5]));
 sky130_fd_sc_hd__buf_4 _3026_ (.A(net449),
    .X(dst_wdata[6]));
 sky130_fd_sc_hd__buf_4 _3027_ (.A(net450),
    .X(dst_wdata[7]));
 sky130_fd_sc_hd__buf_4 _3028_ (.A(net451),
    .X(dst_wdata[8]));
 sky130_fd_sc_hd__buf_4 _3029_ (.A(net452),
    .X(dst_wdata[9]));
 sky130_fd_sc_hd__buf_4 _3030_ (.A(net453),
    .X(dst_wdata[10]));
 sky130_fd_sc_hd__buf_4 _3031_ (.A(net454),
    .X(dst_wdata[11]));
 sky130_fd_sc_hd__buf_4 _3032_ (.A(net455),
    .X(dst_wdata[12]));
 sky130_fd_sc_hd__buf_4 _3033_ (.A(net456),
    .X(dst_wdata[13]));
 sky130_fd_sc_hd__buf_4 _3034_ (.A(net457),
    .X(dst_wdata[14]));
 sky130_fd_sc_hd__buf_4 _3035_ (.A(net458),
    .X(dst_wdata[15]));
 sky130_fd_sc_hd__buf_4 _3036_ (.A(net459),
    .X(dst_wdata[16]));
 sky130_fd_sc_hd__buf_4 _3037_ (.A(net460),
    .X(dst_wdata[17]));
 sky130_fd_sc_hd__buf_4 _3038_ (.A(net461),
    .X(dst_wdata[18]));
 sky130_fd_sc_hd__buf_4 _3039_ (.A(net462),
    .X(dst_wdata[19]));
 sky130_fd_sc_hd__buf_4 _3040_ (.A(net463),
    .X(dst_wdata[20]));
 sky130_fd_sc_hd__buf_4 _3041_ (.A(net464),
    .X(dst_wdata[21]));
 sky130_fd_sc_hd__buf_4 _3042_ (.A(net465),
    .X(dst_wdata[22]));
 sky130_fd_sc_hd__buf_4 _3043_ (.A(net466),
    .X(dst_wdata[23]));
 sky130_fd_sc_hd__buf_4 _3044_ (.A(net467),
    .X(dst_wdata[24]));
 sky130_fd_sc_hd__buf_4 _3045_ (.A(net468),
    .X(dst_wdata[25]));
 sky130_fd_sc_hd__buf_4 _3046_ (.A(net469),
    .X(dst_wdata[26]));
 sky130_fd_sc_hd__buf_4 _3047_ (.A(net470),
    .X(dst_wdata[27]));
 sky130_fd_sc_hd__buf_4 _3048_ (.A(net471),
    .X(dst_wdata[28]));
 sky130_fd_sc_hd__buf_4 _3049_ (.A(net472),
    .X(dst_wdata[29]));
 sky130_fd_sc_hd__buf_4 _3050_ (.A(net473),
    .X(dst_wdata[30]));
 sky130_fd_sc_hd__buf_4 _3051_ (.A(net474),
    .X(dst_wdata[31]));
 sky130_fd_sc_hd__buf_4 _3052_ (.A(net475),
    .X(dst_wdata[32]));
 sky130_fd_sc_hd__buf_4 _3053_ (.A(net476),
    .X(dst_wdata[33]));
 sky130_fd_sc_hd__buf_4 _3054_ (.A(net477),
    .X(dst_wdata[34]));
 sky130_fd_sc_hd__buf_4 _3055_ (.A(net478),
    .X(dst_wdata[35]));
 sky130_fd_sc_hd__buf_4 _3056_ (.A(net479),
    .X(dst_wdata[36]));
 sky130_fd_sc_hd__buf_4 _3057_ (.A(net480),
    .X(dst_wdata[37]));
 sky130_fd_sc_hd__buf_4 _3058_ (.A(net481),
    .X(dst_wdata[38]));
 sky130_fd_sc_hd__buf_4 _3059_ (.A(net482),
    .X(dst_wdata[39]));
 sky130_fd_sc_hd__buf_4 _3060_ (.A(net483),
    .X(dst_wdata[40]));
 sky130_fd_sc_hd__buf_4 _3061_ (.A(net484),
    .X(dst_wdata[41]));
 sky130_fd_sc_hd__buf_4 _3062_ (.A(net485),
    .X(dst_wdata[42]));
 sky130_fd_sc_hd__buf_4 _3063_ (.A(net486),
    .X(dst_wdata[43]));
 sky130_fd_sc_hd__buf_4 _3064_ (.A(net487),
    .X(dst_wdata[44]));
 sky130_fd_sc_hd__buf_4 _3065_ (.A(net488),
    .X(dst_wdata[45]));
 sky130_fd_sc_hd__buf_4 _3066_ (.A(net489),
    .X(dst_wdata[46]));
 sky130_fd_sc_hd__buf_4 _3067_ (.A(net490),
    .X(dst_wdata[47]));
 sky130_fd_sc_hd__buf_4 _3068_ (.A(net491),
    .X(dst_wdata[48]));
 sky130_fd_sc_hd__buf_4 _3069_ (.A(net492),
    .X(dst_wdata[49]));
 sky130_fd_sc_hd__buf_4 _3070_ (.A(net493),
    .X(dst_wdata[50]));
 sky130_fd_sc_hd__buf_4 _3071_ (.A(net494),
    .X(dst_wdata[51]));
 sky130_fd_sc_hd__buf_4 _3072_ (.A(net495),
    .X(dst_wdata[52]));
 sky130_fd_sc_hd__buf_4 _3073_ (.A(net496),
    .X(dst_wdata[53]));
 sky130_fd_sc_hd__buf_4 _3074_ (.A(net497),
    .X(dst_wdata[54]));
 sky130_fd_sc_hd__buf_4 _3075_ (.A(net498),
    .X(dst_wdata[55]));
 sky130_fd_sc_hd__buf_4 _3076_ (.A(net499),
    .X(dst_wdata[56]));
 sky130_fd_sc_hd__buf_4 _3077_ (.A(net500),
    .X(dst_wdata[57]));
 sky130_fd_sc_hd__buf_4 _3078_ (.A(net501),
    .X(dst_wdata[58]));
 sky130_fd_sc_hd__buf_4 _3079_ (.A(net502),
    .X(dst_wdata[59]));
 sky130_fd_sc_hd__buf_4 _3080_ (.A(net503),
    .X(dst_wdata[60]));
 sky130_fd_sc_hd__buf_4 _3081_ (.A(net504),
    .X(dst_wdata[61]));
 sky130_fd_sc_hd__buf_4 _3082_ (.A(net505),
    .X(dst_wdata[62]));
 sky130_fd_sc_hd__buf_4 _3083_ (.A(net506),
    .X(dst_wdata[63]));
 sky130_fd_sc_hd__buf_4 _3084_ (.A(net507),
    .X(dst_wdata[64]));
 sky130_fd_sc_hd__buf_4 _3085_ (.A(net508),
    .X(dst_wdata[65]));
 sky130_fd_sc_hd__buf_4 _3086_ (.A(net509),
    .X(dst_wdata[66]));
 sky130_fd_sc_hd__buf_4 _3087_ (.A(net510),
    .X(dst_wdata[67]));
 sky130_fd_sc_hd__buf_4 _3088_ (.A(net511),
    .X(dst_wdata[68]));
 sky130_fd_sc_hd__buf_4 _3089_ (.A(net512),
    .X(dst_wdata[69]));
 sky130_fd_sc_hd__buf_4 _3090_ (.A(net513),
    .X(dst_wdata[70]));
 sky130_fd_sc_hd__buf_4 _3091_ (.A(net514),
    .X(dst_wdata[71]));
 sky130_fd_sc_hd__buf_4 _3092_ (.A(net515),
    .X(dst_wdata[72]));
 sky130_fd_sc_hd__buf_4 _3093_ (.A(net516),
    .X(dst_wdata[73]));
 sky130_fd_sc_hd__buf_4 _3094_ (.A(net517),
    .X(dst_wdata[74]));
 sky130_fd_sc_hd__buf_4 _3095_ (.A(net518),
    .X(dst_wdata[75]));
 sky130_fd_sc_hd__buf_4 _3096_ (.A(net519),
    .X(dst_wdata[76]));
 sky130_fd_sc_hd__buf_4 _3097_ (.A(net520),
    .X(dst_wdata[77]));
 sky130_fd_sc_hd__buf_4 _3098_ (.A(net521),
    .X(dst_wdata[78]));
 sky130_fd_sc_hd__buf_4 _3099_ (.A(net522),
    .X(dst_wdata[79]));
 sky130_fd_sc_hd__buf_4 _3100_ (.A(net523),
    .X(dst_wdata[80]));
 sky130_fd_sc_hd__buf_4 _3101_ (.A(net524),
    .X(dst_wdata[81]));
 sky130_fd_sc_hd__buf_4 _3102_ (.A(net525),
    .X(dst_wdata[82]));
 sky130_fd_sc_hd__buf_4 _3103_ (.A(net526),
    .X(dst_wdata[83]));
 sky130_fd_sc_hd__buf_4 _3104_ (.A(net527),
    .X(dst_wdata[84]));
 sky130_fd_sc_hd__buf_4 _3105_ (.A(net528),
    .X(dst_wdata[85]));
 sky130_fd_sc_hd__buf_4 _3106_ (.A(net529),
    .X(dst_wdata[86]));
 sky130_fd_sc_hd__buf_4 _3107_ (.A(net530),
    .X(dst_wdata[87]));
 sky130_fd_sc_hd__buf_4 _3108_ (.A(net531),
    .X(dst_wdata[88]));
 sky130_fd_sc_hd__buf_4 _3109_ (.A(net532),
    .X(dst_wdata[89]));
 sky130_fd_sc_hd__buf_4 _3110_ (.A(net533),
    .X(dst_wdata[90]));
 sky130_fd_sc_hd__buf_4 _3111_ (.A(net534),
    .X(dst_wdata[91]));
 sky130_fd_sc_hd__buf_4 _3112_ (.A(net535),
    .X(dst_wdata[92]));
 sky130_fd_sc_hd__buf_4 _3113_ (.A(net536),
    .X(dst_wdata[93]));
 sky130_fd_sc_hd__buf_4 _3114_ (.A(net537),
    .X(dst_wdata[94]));
 sky130_fd_sc_hd__buf_4 _3115_ (.A(net538),
    .X(dst_wdata[95]));
 sky130_fd_sc_hd__buf_4 _3116_ (.A(net539),
    .X(dst_wdata[96]));
 sky130_fd_sc_hd__buf_4 _3117_ (.A(net540),
    .X(dst_wdata[97]));
 sky130_fd_sc_hd__buf_4 _3118_ (.A(net541),
    .X(dst_wdata[98]));
 sky130_fd_sc_hd__buf_4 _3119_ (.A(net542),
    .X(dst_wdata[99]));
 sky130_fd_sc_hd__buf_4 _3120_ (.A(net543),
    .X(dst_wdata[100]));
 sky130_fd_sc_hd__buf_4 _3121_ (.A(net544),
    .X(dst_wdata[101]));
 sky130_fd_sc_hd__buf_4 _3122_ (.A(net545),
    .X(dst_wdata[102]));
 sky130_fd_sc_hd__buf_4 _3123_ (.A(net546),
    .X(dst_wdata[103]));
 sky130_fd_sc_hd__buf_4 _3124_ (.A(net547),
    .X(dst_wdata[104]));
 sky130_fd_sc_hd__buf_4 _3125_ (.A(net548),
    .X(dst_wdata[105]));
 sky130_fd_sc_hd__buf_4 _3126_ (.A(net549),
    .X(dst_wdata[106]));
 sky130_fd_sc_hd__buf_4 _3127_ (.A(net550),
    .X(dst_wdata[107]));
 sky130_fd_sc_hd__buf_4 _3128_ (.A(net551),
    .X(dst_wdata[108]));
 sky130_fd_sc_hd__buf_4 _3129_ (.A(net552),
    .X(dst_wdata[109]));
 sky130_fd_sc_hd__buf_4 _3130_ (.A(net553),
    .X(dst_wdata[110]));
 sky130_fd_sc_hd__buf_4 _3131_ (.A(net554),
    .X(dst_wdata[111]));
 sky130_fd_sc_hd__buf_4 _3132_ (.A(net555),
    .X(dst_wdata[112]));
 sky130_fd_sc_hd__buf_4 _3133_ (.A(net556),
    .X(dst_wdata[113]));
 sky130_fd_sc_hd__buf_4 _3134_ (.A(net557),
    .X(dst_wdata[114]));
 sky130_fd_sc_hd__buf_4 _3135_ (.A(net558),
    .X(dst_wdata[115]));
 sky130_fd_sc_hd__buf_4 _3136_ (.A(net559),
    .X(dst_wdata[116]));
 sky130_fd_sc_hd__buf_4 _3137_ (.A(net560),
    .X(dst_wdata[117]));
 sky130_fd_sc_hd__buf_4 _3138_ (.A(net561),
    .X(dst_wdata[118]));
 sky130_fd_sc_hd__buf_4 _3139_ (.A(net562),
    .X(dst_wdata[119]));
 sky130_fd_sc_hd__buf_4 _3140_ (.A(net563),
    .X(dst_wdata[120]));
 sky130_fd_sc_hd__buf_4 _3141_ (.A(net564),
    .X(dst_wdata[121]));
 sky130_fd_sc_hd__buf_4 _3142_ (.A(net565),
    .X(dst_wdata[122]));
 sky130_fd_sc_hd__buf_4 _3143_ (.A(net566),
    .X(dst_wdata[123]));
 sky130_fd_sc_hd__buf_4 _3144_ (.A(net567),
    .X(dst_wdata[124]));
 sky130_fd_sc_hd__buf_4 _3145_ (.A(net568),
    .X(dst_wdata[125]));
 sky130_fd_sc_hd__buf_4 _3146_ (.A(net569),
    .X(dst_wdata[126]));
 sky130_fd_sc_hd__buf_4 _3147_ (.A(net570),
    .X(dst_wdata[127]));
 sky130_fd_sc_hd__buf_4 _3148_ (.A(net571),
    .X(dst_wstrb[0]));
 sky130_fd_sc_hd__buf_4 _3149_ (.A(net572),
    .X(dst_wstrb[1]));
 sky130_fd_sc_hd__buf_4 _3150_ (.A(net573),
    .X(dst_wstrb[2]));
 sky130_fd_sc_hd__buf_4 _3151_ (.A(net574),
    .X(dst_wstrb[3]));
 sky130_fd_sc_hd__buf_4 _3152_ (.A(net575),
    .X(dst_wstrb[4]));
 sky130_fd_sc_hd__buf_4 _3153_ (.A(net576),
    .X(dst_wstrb[5]));
 sky130_fd_sc_hd__buf_4 _3154_ (.A(net577),
    .X(dst_wstrb[6]));
 sky130_fd_sc_hd__buf_4 _3155_ (.A(net578),
    .X(dst_wstrb[7]));
 sky130_fd_sc_hd__buf_4 _3156_ (.A(net579),
    .X(dst_wstrb[8]));
 sky130_fd_sc_hd__buf_4 _3157_ (.A(net580),
    .X(dst_wstrb[9]));
 sky130_fd_sc_hd__buf_4 _3158_ (.A(net581),
    .X(dst_wstrb[10]));
 sky130_fd_sc_hd__buf_4 _3159_ (.A(net582),
    .X(dst_wstrb[11]));
 sky130_fd_sc_hd__buf_4 _3160_ (.A(net583),
    .X(dst_wstrb[12]));
 sky130_fd_sc_hd__buf_4 _3161_ (.A(net584),
    .X(dst_wstrb[13]));
 sky130_fd_sc_hd__buf_4 _3162_ (.A(net585),
    .X(dst_wstrb[14]));
 sky130_fd_sc_hd__buf_4 _3163_ (.A(net586),
    .X(dst_wstrb[15]));
 sky130_fd_sc_hd__buf_4 _3164_ (.A(net587),
    .X(src_addr[0]));
 sky130_fd_sc_hd__buf_4 _3165_ (.A(net588),
    .X(src_addr[1]));
 sky130_fd_sc_hd__buf_4 _3166_ (.A(net589),
    .X(src_addr[2]));
 sky130_fd_sc_hd__buf_4 _3167_ (.A(net590),
    .X(src_addr[3]));
 sky130_fd_sc_hd__buf_4 _3168_ (.A(net591),
    .X(src_addr[4]));
 sky130_fd_sc_hd__buf_4 _3169_ (.A(net592),
    .X(src_addr[5]));
 sky130_fd_sc_hd__buf_4 _3170_ (.A(net593),
    .X(src_addr[6]));
 sky130_fd_sc_hd__buf_4 _3171_ (.A(net594),
    .X(src_addr[7]));
 sky130_fd_sc_hd__buf_4 _3172_ (.A(net595),
    .X(src_addr[8]));
 sky130_fd_sc_hd__buf_4 _3173_ (.A(net596),
    .X(src_addr[9]));
 sky130_fd_sc_hd__buf_4 _3174_ (.A(net597),
    .X(src_addr[10]));
 sky130_fd_sc_hd__buf_4 _3175_ (.A(net598),
    .X(src_addr[11]));
 sky130_fd_sc_hd__buf_4 _3176_ (.A(net599),
    .X(src_addr[12]));
 sky130_fd_sc_hd__buf_4 _3177_ (.A(net600),
    .X(src_addr[13]));
 sky130_fd_sc_hd__buf_4 _3178_ (.A(net601),
    .X(src_addr[14]));
 sky130_fd_sc_hd__buf_4 _3179_ (.A(net602),
    .X(src_addr[15]));
 sky130_fd_sc_hd__buf_4 _3180_ (.A(net603),
    .X(src_addr[16]));
 sky130_fd_sc_hd__buf_4 _3181_ (.A(net604),
    .X(src_addr[17]));
 sky130_fd_sc_hd__buf_4 _3182_ (.A(net605),
    .X(src_addr[18]));
 sky130_fd_sc_hd__buf_4 _3183_ (.A(net606),
    .X(src_addr[19]));
 sky130_fd_sc_hd__buf_4 _3184_ (.A(net607),
    .X(src_addr[20]));
 sky130_fd_sc_hd__buf_4 _3185_ (.A(net608),
    .X(src_addr[21]));
 sky130_fd_sc_hd__buf_4 _3186_ (.A(net609),
    .X(src_addr[22]));
 sky130_fd_sc_hd__buf_4 _3187_ (.A(net610),
    .X(src_addr[23]));
 sky130_fd_sc_hd__buf_4 _3188_ (.A(net611),
    .X(src_addr[24]));
 sky130_fd_sc_hd__buf_4 _3189_ (.A(net612),
    .X(src_addr[25]));
 sky130_fd_sc_hd__buf_4 _3190_ (.A(net613),
    .X(src_addr[26]));
 sky130_fd_sc_hd__buf_4 _3191_ (.A(net614),
    .X(src_addr[27]));
 sky130_fd_sc_hd__buf_4 _3192_ (.A(net615),
    .X(src_addr[28]));
 sky130_fd_sc_hd__buf_4 _3193_ (.A(net616),
    .X(src_addr[29]));
 sky130_fd_sc_hd__buf_4 _3194_ (.A(net617),
    .X(src_addr[30]));
 sky130_fd_sc_hd__buf_4 _3195_ (.A(net618),
    .X(src_addr[31]));
 sky130_fd_sc_hd__buf_4 _3196_ (.A(net619),
    .X(src_addr[32]));
 sky130_fd_sc_hd__buf_4 _3197_ (.A(net620),
    .X(src_addr[33]));
 sky130_fd_sc_hd__buf_4 _3198_ (.A(net621),
    .X(src_addr[34]));
 sky130_fd_sc_hd__buf_4 _3199_ (.A(net622),
    .X(src_addr[35]));
 sky130_fd_sc_hd__buf_4 _3200_ (.A(net623),
    .X(src_addr[36]));
 sky130_fd_sc_hd__buf_4 _3201_ (.A(net624),
    .X(src_addr[37]));
 sky130_fd_sc_hd__buf_4 _3202_ (.A(net625),
    .X(src_addr[38]));
 sky130_fd_sc_hd__buf_4 _3203_ (.A(net626),
    .X(src_addr[39]));
 sky130_fd_sc_hd__buf_4 _3204_ (.A(net627),
    .X(src_addr[40]));
 sky130_fd_sc_hd__buf_4 _3205_ (.A(net628),
    .X(src_addr[41]));
 sky130_fd_sc_hd__buf_4 _3206_ (.A(net629),
    .X(src_addr[42]));
 sky130_fd_sc_hd__buf_4 _3207_ (.A(net630),
    .X(src_addr[43]));
 sky130_fd_sc_hd__buf_4 _3208_ (.A(net631),
    .X(src_addr[44]));
 sky130_fd_sc_hd__buf_4 _3209_ (.A(net632),
    .X(src_addr[45]));
 sky130_fd_sc_hd__buf_4 _3210_ (.A(net633),
    .X(src_addr[46]));
 sky130_fd_sc_hd__buf_4 _3211_ (.A(net634),
    .X(src_addr[47]));
 sky130_fd_sc_hd__buf_4 _3212_ (.A(net635),
    .X(src_addr[48]));
 sky130_fd_sc_hd__buf_4 _3213_ (.A(net636),
    .X(src_addr[49]));
 sky130_fd_sc_hd__buf_4 _3214_ (.A(net637),
    .X(src_addr[50]));
 sky130_fd_sc_hd__buf_4 _3215_ (.A(net638),
    .X(src_addr[51]));
 sky130_fd_sc_hd__buf_4 _3216_ (.A(net639),
    .X(src_addr[52]));
 sky130_fd_sc_hd__buf_4 _3217_ (.A(net640),
    .X(src_addr[53]));
 sky130_fd_sc_hd__buf_4 _3218_ (.A(net641),
    .X(src_addr[54]));
 sky130_fd_sc_hd__buf_4 _3219_ (.A(net642),
    .X(src_addr[55]));
 sky130_fd_sc_hd__buf_4 _3220_ (.A(net643),
    .X(src_addr[56]));
 sky130_fd_sc_hd__buf_4 _3221_ (.A(net644),
    .X(src_addr[57]));
 sky130_fd_sc_hd__buf_4 _3222_ (.A(net645),
    .X(src_addr[58]));
 sky130_fd_sc_hd__buf_4 _3223_ (.A(net646),
    .X(src_addr[59]));
 sky130_fd_sc_hd__buf_4 _3224_ (.A(net647),
    .X(src_addr[60]));
 sky130_fd_sc_hd__buf_4 _3225_ (.A(net648),
    .X(src_addr[61]));
 sky130_fd_sc_hd__buf_4 _3226_ (.A(net649),
    .X(src_addr[62]));
 sky130_fd_sc_hd__buf_4 _3227_ (.A(net650),
    .X(src_addr[63]));
 sky130_fd_sc_hd__buf_4 _3228_ (.A(net651),
    .X(src_addr[64]));
 sky130_fd_sc_hd__buf_4 _3229_ (.A(net652),
    .X(src_addr[65]));
 sky130_fd_sc_hd__buf_4 _3230_ (.A(net653),
    .X(src_addr[66]));
 sky130_fd_sc_hd__buf_4 _3231_ (.A(net654),
    .X(src_addr[67]));
 sky130_fd_sc_hd__buf_4 _3232_ (.A(net655),
    .X(src_addr[68]));
 sky130_fd_sc_hd__buf_4 _3233_ (.A(net656),
    .X(src_addr[69]));
 sky130_fd_sc_hd__buf_4 _3234_ (.A(net657),
    .X(src_addr[70]));
 sky130_fd_sc_hd__buf_4 _3235_ (.A(net658),
    .X(src_addr[71]));
 sky130_fd_sc_hd__buf_4 _3236_ (.A(net659),
    .X(src_addr[72]));
 sky130_fd_sc_hd__buf_4 _3237_ (.A(net660),
    .X(src_addr[73]));
 sky130_fd_sc_hd__buf_4 _3238_ (.A(net661),
    .X(src_addr[74]));
 sky130_fd_sc_hd__buf_4 _3239_ (.A(net662),
    .X(src_addr[75]));
 sky130_fd_sc_hd__buf_4 _3240_ (.A(net663),
    .X(src_addr[76]));
 sky130_fd_sc_hd__buf_4 _3241_ (.A(net664),
    .X(src_addr[77]));
 sky130_fd_sc_hd__buf_4 _3242_ (.A(net665),
    .X(src_addr[78]));
 sky130_fd_sc_hd__buf_4 _3243_ (.A(net666),
    .X(src_addr[79]));
 sky130_fd_sc_hd__buf_4 _3244_ (.A(net667),
    .X(src_addr[80]));
 sky130_fd_sc_hd__buf_4 _3245_ (.A(net668),
    .X(src_addr[81]));
 sky130_fd_sc_hd__buf_4 _3246_ (.A(net669),
    .X(src_addr[82]));
 sky130_fd_sc_hd__buf_4 _3247_ (.A(net670),
    .X(src_addr[83]));
 sky130_fd_sc_hd__buf_4 _3248_ (.A(net671),
    .X(src_addr[84]));
 sky130_fd_sc_hd__buf_4 _3249_ (.A(net672),
    .X(src_addr[85]));
 sky130_fd_sc_hd__buf_4 _3250_ (.A(net673),
    .X(src_addr[86]));
 sky130_fd_sc_hd__buf_4 _3251_ (.A(net674),
    .X(src_addr[87]));
 sky130_fd_sc_hd__buf_4 _3252_ (.A(net675),
    .X(src_addr[88]));
 sky130_fd_sc_hd__buf_4 _3253_ (.A(net676),
    .X(src_addr[89]));
 sky130_fd_sc_hd__buf_4 _3254_ (.A(net677),
    .X(src_addr[90]));
 sky130_fd_sc_hd__buf_4 _3255_ (.A(net678),
    .X(src_addr[91]));
 sky130_fd_sc_hd__buf_4 _3256_ (.A(net679),
    .X(src_addr[92]));
 sky130_fd_sc_hd__buf_4 _3257_ (.A(net680),
    .X(src_addr[93]));
 sky130_fd_sc_hd__buf_4 _3258_ (.A(net681),
    .X(src_addr[94]));
 sky130_fd_sc_hd__buf_4 _3259_ (.A(net682),
    .X(src_addr[95]));
 sky130_fd_sc_hd__buf_4 _3260_ (.A(net683),
    .X(src_addr[96]));
 sky130_fd_sc_hd__buf_4 _3261_ (.A(net684),
    .X(src_addr[97]));
 sky130_fd_sc_hd__buf_4 _3262_ (.A(net685),
    .X(src_addr[98]));
 sky130_fd_sc_hd__buf_4 _3263_ (.A(net686),
    .X(src_addr[99]));
 sky130_fd_sc_hd__buf_4 _3264_ (.A(net687),
    .X(src_addr[100]));
 sky130_fd_sc_hd__buf_4 _3265_ (.A(net688),
    .X(src_addr[101]));
 sky130_fd_sc_hd__buf_4 _3266_ (.A(net689),
    .X(src_addr[102]));
 sky130_fd_sc_hd__buf_4 _3267_ (.A(net690),
    .X(src_addr[103]));
 sky130_fd_sc_hd__buf_4 _3268_ (.A(net691),
    .X(src_addr[104]));
 sky130_fd_sc_hd__buf_4 _3269_ (.A(net692),
    .X(src_addr[105]));
 sky130_fd_sc_hd__buf_4 _3270_ (.A(net693),
    .X(src_addr[106]));
 sky130_fd_sc_hd__buf_4 _3271_ (.A(net694),
    .X(src_addr[107]));
 sky130_fd_sc_hd__buf_4 _3272_ (.A(net695),
    .X(src_addr[108]));
 sky130_fd_sc_hd__buf_4 _3273_ (.A(net696),
    .X(src_addr[109]));
 sky130_fd_sc_hd__buf_4 _3274_ (.A(net697),
    .X(src_addr[110]));
 sky130_fd_sc_hd__buf_4 _3275_ (.A(net698),
    .X(src_addr[111]));
 sky130_fd_sc_hd__buf_4 _3276_ (.A(net699),
    .X(src_addr[112]));
 sky130_fd_sc_hd__buf_4 _3277_ (.A(net700),
    .X(src_addr[113]));
 sky130_fd_sc_hd__buf_4 _3278_ (.A(net701),
    .X(src_addr[114]));
 sky130_fd_sc_hd__buf_4 _3279_ (.A(net702),
    .X(src_addr[115]));
 sky130_fd_sc_hd__buf_4 _3280_ (.A(net703),
    .X(src_addr[116]));
 sky130_fd_sc_hd__buf_4 _3281_ (.A(net704),
    .X(src_addr[117]));
 sky130_fd_sc_hd__buf_4 _3282_ (.A(net705),
    .X(src_addr[118]));
 sky130_fd_sc_hd__buf_4 _3283_ (.A(net706),
    .X(src_addr[119]));
 sky130_fd_sc_hd__buf_4 _3284_ (.A(net707),
    .X(src_addr[120]));
 sky130_fd_sc_hd__buf_4 _3285_ (.A(net708),
    .X(src_addr[121]));
 sky130_fd_sc_hd__buf_4 _3286_ (.A(net709),
    .X(src_addr[122]));
 sky130_fd_sc_hd__buf_4 _3287_ (.A(net710),
    .X(src_addr[123]));
 sky130_fd_sc_hd__buf_4 _3288_ (.A(net711),
    .X(src_addr[124]));
 sky130_fd_sc_hd__buf_4 _3289_ (.A(net712),
    .X(src_addr[125]));
 sky130_fd_sc_hd__buf_4 _3290_ (.A(net713),
    .X(src_addr[126]));
 sky130_fd_sc_hd__buf_4 _3291_ (.A(net714),
    .X(src_addr[127]));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[0]$_DFF_PN0_  (.D(_0000_),
    .Q(\active_channel_count[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[1]$_DFF_PN0_  (.D(_0001_),
    .Q(\active_channel_count[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[2]$_DFF_PN0_  (.D(_0002_),
    .Q(\active_channel_count[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[3]$_DFF_PN0_  (.D(_0003_),
    .Q(\active_channel_count[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[0]$_DFF_PN0_  (.D(_0004_),
    .Q(net146),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[1]$_DFF_PN0_  (.D(_0005_),
    .Q(net147),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[2]$_DFF_PN0_  (.D(_0006_),
    .Q(net148),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \channel_busy[3]$_DFF_PN0_  (.D(_0007_),
    .Q(net149),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[0]$_DFF_PN0_  (.D(_1441_),
    .Q(net150),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[1]$_DFF_PN0_  (.D(_1439_),
    .Q(net151),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[2]$_DFF_PN0_  (.D(_1436_),
    .Q(net152),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[3]$_DFF_PN0_  (.D(_1438_),
    .Q(net153),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[0]$_DFF_PN0_  (.D(_0008_),
    .Q(net154),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[1]$_DFF_PN0_  (.D(_0009_),
    .Q(net155),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[2]$_DFF_PN0_  (.D(_0010_),
    .Q(net156),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \channel_error[3]$_DFF_PN0_  (.D(_0011_),
    .Q(net157),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][0]$_DFF_PN0_  (.D(_1030_),
    .Q(\channel_state[0][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][1]$_DFF_PN0_  (.D(_1031_),
    .Q(\channel_state[0][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][2]$_DFF_PN0_  (.D(_1032_),
    .Q(\channel_state[0][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][0]$_DFF_PN0_  (.D(_1027_),
    .Q(\channel_state[1][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][1]$_DFF_PN0_  (.D(_1028_),
    .Q(\channel_state[1][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][2]$_DFF_PN0_  (.D(_1029_),
    .Q(\channel_state[1][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \channel_state[2][0]$_DFF_PN0_  (.D(_1024_),
    .Q(\channel_state[2][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[2][1]$_DFF_PN0_  (.D(_1025_),
    .Q(\channel_state[2][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[2][2]$_DFF_PN0_  (.D(_1026_),
    .Q(\channel_state[2][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[3][0]$_DFF_PN0_  (.D(_1021_),
    .Q(\channel_state[3][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \channel_state[3][1]$_DFF_PN0_  (.D(_1022_),
    .Q(\channel_state[3][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[3][2]$_DFF_PN0_  (.D(_1023_),
    .Q(\channel_state[3][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[0]$_DFF_PN0_  (.D(\active_channel_count[0] ),
    .Q(net158),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[1]$_DFF_PN0_  (.D(\active_channel_count[1] ),
    .Q(net159),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[2]$_DFF_PN0_  (.D(\active_channel_count[2] ),
    .Q(net160),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[3]$_DFF_PN0_  (.D(\active_channel_count[3] ),
    .Q(net161),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_has_active_channels$_DFF_PN0_  (.D(_0012_),
    .Q(net162),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[0]$_DFFE_PN0P_  (.D(_0141_),
    .Q(net163),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[1]$_DFFE_PN0P_  (.D(_0142_),
    .Q(net164),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[2]$_DFFE_PN0P_  (.D(_0143_),
    .Q(net165),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \dst_write[3]$_DFFE_PN0P_  (.D(_0144_),
    .Q(net166),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \src_read[0]$_DFF_PN0_  (.D(_1019_),
    .Q(net167),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_read[1]$_DFF_PN0_  (.D(_1018_),
    .Q(net168),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_read[2]$_DFF_PN0_  (.D(_1017_),
    .Q(net169),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_read[3]$_DFF_PN0_  (.D(_1020_),
    .Q(net170),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \src_rready[0]$_DFF_PN0_  (.D(_1442_),
    .Q(net171),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_rready[1]$_DFF_PN0_  (.D(_1440_),
    .Q(net172),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_rready[2]$_DFF_PN0_  (.D(_1437_),
    .Q(net173),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \src_rready[3]$_DFFE_PN0P_  (.D(_0145_),
    .Q(net174),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][0]$_DFF_PN0_  (.D(_0013_),
    .Q(\transfer_count[0][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][10]$_DFF_PN0_  (.D(_0014_),
    .Q(\transfer_count[0][10] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][11]$_DFF_PN0_  (.D(_0015_),
    .Q(\transfer_count[0][11] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][12]$_DFF_PN0_  (.D(_0016_),
    .Q(\transfer_count[0][12] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][13]$_DFF_PN0_  (.D(_0017_),
    .Q(\transfer_count[0][13] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][14]$_DFF_PN0_  (.D(_0018_),
    .Q(\transfer_count[0][14] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][15]$_DFF_PN0_  (.D(_0019_),
    .Q(\transfer_count[0][15] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][16]$_DFF_PN0_  (.D(_0020_),
    .Q(\transfer_count[0][16] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][17]$_DFF_PN0_  (.D(_0021_),
    .Q(\transfer_count[0][17] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][18]$_DFF_PN0_  (.D(_0022_),
    .Q(\transfer_count[0][18] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][19]$_DFF_PN0_  (.D(_0023_),
    .Q(\transfer_count[0][19] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][1]$_DFF_PN0_  (.D(_0024_),
    .Q(\transfer_count[0][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][20]$_DFF_PN0_  (.D(_0025_),
    .Q(\transfer_count[0][20] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][21]$_DFF_PN0_  (.D(_0026_),
    .Q(\transfer_count[0][21] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][22]$_DFF_PN0_  (.D(_0027_),
    .Q(\transfer_count[0][22] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][23]$_DFF_PN0_  (.D(_0028_),
    .Q(\transfer_count[0][23] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][24]$_DFF_PN0_  (.D(_0029_),
    .Q(\transfer_count[0][24] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][25]$_DFF_PN0_  (.D(_0030_),
    .Q(\transfer_count[0][25] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][26]$_DFF_PN0_  (.D(_0031_),
    .Q(\transfer_count[0][26] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][27]$_DFF_PN0_  (.D(_0032_),
    .Q(\transfer_count[0][27] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][28]$_DFF_PN0_  (.D(_0033_),
    .Q(\transfer_count[0][28] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][29]$_DFF_PN0_  (.D(_0034_),
    .Q(\transfer_count[0][29] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \transfer_count[0][2]$_DFF_PN0_  (.D(_0035_),
    .Q(\transfer_count[0][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][30]$_DFF_PN0_  (.D(_0036_),
    .Q(\transfer_count[0][30] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][31]$_DFF_PN0_  (.D(_0037_),
    .Q(\transfer_count[0][31] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][3]$_DFF_PN0_  (.D(_0038_),
    .Q(\transfer_count[0][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][4]$_DFF_PN0_  (.D(_0039_),
    .Q(\transfer_count[0][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][5]$_DFF_PN0_  (.D(_0040_),
    .Q(\transfer_count[0][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[0][6]$_DFF_PN0_  (.D(_0041_),
    .Q(\transfer_count[0][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][7]$_DFF_PN0_  (.D(_0042_),
    .Q(\transfer_count[0][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][8]$_DFF_PN0_  (.D(_0043_),
    .Q(\transfer_count[0][8] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][9]$_DFF_PN0_  (.D(_0044_),
    .Q(\transfer_count[0][9] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][0]$_DFF_PN0_  (.D(_0045_),
    .Q(\transfer_count[1][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][10]$_DFF_PN0_  (.D(_0046_),
    .Q(\transfer_count[1][10] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][11]$_DFF_PN0_  (.D(_0047_),
    .Q(\transfer_count[1][11] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][12]$_DFF_PN0_  (.D(_0048_),
    .Q(\transfer_count[1][12] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][13]$_DFF_PN0_  (.D(_0049_),
    .Q(\transfer_count[1][13] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][14]$_DFF_PN0_  (.D(_0050_),
    .Q(\transfer_count[1][14] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][15]$_DFF_PN0_  (.D(_0051_),
    .Q(\transfer_count[1][15] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][16]$_DFF_PN0_  (.D(_0052_),
    .Q(\transfer_count[1][16] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][17]$_DFF_PN0_  (.D(_0053_),
    .Q(\transfer_count[1][17] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[1][18]$_DFF_PN0_  (.D(_0054_),
    .Q(\transfer_count[1][18] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][19]$_DFF_PN0_  (.D(_0055_),
    .Q(\transfer_count[1][19] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][1]$_DFF_PN0_  (.D(_0056_),
    .Q(\transfer_count[1][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][20]$_DFF_PN0_  (.D(_0057_),
    .Q(\transfer_count[1][20] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][21]$_DFF_PN0_  (.D(_0058_),
    .Q(\transfer_count[1][21] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][22]$_DFF_PN0_  (.D(_0059_),
    .Q(\transfer_count[1][22] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[1][23]$_DFF_PN0_  (.D(_0060_),
    .Q(\transfer_count[1][23] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][24]$_DFF_PN0_  (.D(_0061_),
    .Q(\transfer_count[1][24] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][25]$_DFF_PN0_  (.D(_0062_),
    .Q(\transfer_count[1][25] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][26]$_DFF_PN0_  (.D(_0063_),
    .Q(\transfer_count[1][26] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][27]$_DFF_PN0_  (.D(_0064_),
    .Q(\transfer_count[1][27] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][28]$_DFF_PN0_  (.D(_0065_),
    .Q(\transfer_count[1][28] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][29]$_DFF_PN0_  (.D(_0066_),
    .Q(\transfer_count[1][29] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[1][2]$_DFF_PN0_  (.D(_0067_),
    .Q(\transfer_count[1][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][30]$_DFF_PN0_  (.D(_0068_),
    .Q(\transfer_count[1][30] ),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][31]$_DFF_PN0_  (.D(_0069_),
    .Q(\transfer_count[1][31] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[1][3]$_DFF_PN0_  (.D(_0070_),
    .Q(\transfer_count[1][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][4]$_DFF_PN0_  (.D(_0071_),
    .Q(\transfer_count[1][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][5]$_DFF_PN0_  (.D(_0072_),
    .Q(\transfer_count[1][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][6]$_DFF_PN0_  (.D(_0073_),
    .Q(\transfer_count[1][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][7]$_DFF_PN0_  (.D(_0074_),
    .Q(\transfer_count[1][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[1][8]$_DFF_PN0_  (.D(_0075_),
    .Q(\transfer_count[1][8] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][9]$_DFF_PN0_  (.D(_0076_),
    .Q(\transfer_count[1][9] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][0]$_DFF_PN0_  (.D(_0077_),
    .Q(\transfer_count[2][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][10]$_DFF_PN0_  (.D(_0078_),
    .Q(\transfer_count[2][10] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[2][11]$_DFF_PN0_  (.D(_0079_),
    .Q(\transfer_count[2][11] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][12]$_DFF_PN0_  (.D(_0080_),
    .Q(\transfer_count[2][12] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][13]$_DFF_PN0_  (.D(_0081_),
    .Q(\transfer_count[2][13] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][14]$_DFF_PN0_  (.D(_0082_),
    .Q(\transfer_count[2][14] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][15]$_DFF_PN0_  (.D(_0083_),
    .Q(\transfer_count[2][15] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][16]$_DFF_PN0_  (.D(_0084_),
    .Q(\transfer_count[2][16] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][17]$_DFF_PN0_  (.D(_0085_),
    .Q(\transfer_count[2][17] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][18]$_DFF_PN0_  (.D(_0086_),
    .Q(\transfer_count[2][18] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][19]$_DFF_PN0_  (.D(_0087_),
    .Q(\transfer_count[2][19] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][1]$_DFF_PN0_  (.D(_0088_),
    .Q(\transfer_count[2][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][20]$_DFF_PN0_  (.D(_0089_),
    .Q(\transfer_count[2][20] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][21]$_DFF_PN0_  (.D(_0090_),
    .Q(\transfer_count[2][21] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][22]$_DFF_PN0_  (.D(_0091_),
    .Q(\transfer_count[2][22] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][23]$_DFF_PN0_  (.D(_0092_),
    .Q(\transfer_count[2][23] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][24]$_DFF_PN0_  (.D(_0093_),
    .Q(\transfer_count[2][24] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][25]$_DFF_PN0_  (.D(_0094_),
    .Q(\transfer_count[2][25] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][26]$_DFF_PN0_  (.D(_0095_),
    .Q(\transfer_count[2][26] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][27]$_DFF_PN0_  (.D(_0096_),
    .Q(\transfer_count[2][27] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][28]$_DFF_PN0_  (.D(_0097_),
    .Q(\transfer_count[2][28] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][29]$_DFF_PN0_  (.D(_0098_),
    .Q(\transfer_count[2][29] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][2]$_DFF_PN0_  (.D(_0099_),
    .Q(\transfer_count[2][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][30]$_DFF_PN0_  (.D(_0100_),
    .Q(\transfer_count[2][30] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][31]$_DFF_PN0_  (.D(_0101_),
    .Q(\transfer_count[2][31] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][3]$_DFF_PN0_  (.D(_0102_),
    .Q(\transfer_count[2][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][4]$_DFF_PN0_  (.D(_0103_),
    .Q(\transfer_count[2][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][5]$_DFF_PN0_  (.D(_0104_),
    .Q(\transfer_count[2][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][6]$_DFF_PN0_  (.D(_0105_),
    .Q(\transfer_count[2][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][7]$_DFF_PN0_  (.D(_0106_),
    .Q(\transfer_count[2][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[2][8]$_DFF_PN0_  (.D(_0107_),
    .Q(\transfer_count[2][8] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][9]$_DFF_PN0_  (.D(_0108_),
    .Q(\transfer_count[2][9] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][0]$_DFF_PN0_  (.D(_0109_),
    .Q(\transfer_count[3][0] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][10]$_DFF_PN0_  (.D(_0110_),
    .Q(\transfer_count[3][10] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][11]$_DFF_PN0_  (.D(_0111_),
    .Q(\transfer_count[3][11] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][12]$_DFF_PN0_  (.D(_0112_),
    .Q(\transfer_count[3][12] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][13]$_DFF_PN0_  (.D(_0113_),
    .Q(\transfer_count[3][13] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][14]$_DFF_PN0_  (.D(_0114_),
    .Q(\transfer_count[3][14] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][15]$_DFF_PN0_  (.D(_0115_),
    .Q(\transfer_count[3][15] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][16]$_DFF_PN0_  (.D(_0116_),
    .Q(\transfer_count[3][16] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][17]$_DFF_PN0_  (.D(_0117_),
    .Q(\transfer_count[3][17] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][18]$_DFF_PN0_  (.D(_0118_),
    .Q(\transfer_count[3][18] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][19]$_DFF_PN0_  (.D(_0119_),
    .Q(\transfer_count[3][19] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][1]$_DFF_PN0_  (.D(_0120_),
    .Q(\transfer_count[3][1] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][20]$_DFF_PN0_  (.D(_0121_),
    .Q(\transfer_count[3][20] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][21]$_DFF_PN0_  (.D(_0122_),
    .Q(\transfer_count[3][21] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][22]$_DFF_PN0_  (.D(_0123_),
    .Q(\transfer_count[3][22] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][23]$_DFF_PN0_  (.D(_0124_),
    .Q(\transfer_count[3][23] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][24]$_DFF_PN0_  (.D(_0125_),
    .Q(\transfer_count[3][24] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][25]$_DFF_PN0_  (.D(_0126_),
    .Q(\transfer_count[3][25] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][26]$_DFF_PN0_  (.D(_0127_),
    .Q(\transfer_count[3][26] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][27]$_DFF_PN0_  (.D(_0128_),
    .Q(\transfer_count[3][27] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][28]$_DFF_PN0_  (.D(_0129_),
    .Q(\transfer_count[3][28] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][29]$_DFF_PN0_  (.D(_0130_),
    .Q(\transfer_count[3][29] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \transfer_count[3][2]$_DFF_PN0_  (.D(_0131_),
    .Q(\transfer_count[3][2] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][30]$_DFF_PN0_  (.D(_0132_),
    .Q(\transfer_count[3][30] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][31]$_DFF_PN0_  (.D(_0133_),
    .Q(\transfer_count[3][31] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][3]$_DFF_PN0_  (.D(_0134_),
    .Q(\transfer_count[3][3] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][4]$_DFF_PN0_  (.D(_0135_),
    .Q(\transfer_count[3][4] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][5]$_DFF_PN0_  (.D(_0136_),
    .Q(\transfer_count[3][5] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][6]$_DFF_PN0_  (.D(_0137_),
    .Q(\transfer_count[3][6] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][7]$_DFF_PN0_  (.D(_0138_),
    .Q(\transfer_count[3][7] ),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \transfer_count[3][8]$_DFF_PN0_  (.D(_0139_),
    .Q(\transfer_count[3][8] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][9]$_DFF_PN0_  (.D(_0140_),
    .Q(\transfer_count[3][9] ),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2203 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(channel_enable[0]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(channel_enable[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(channel_enable[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(channel_enable[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(channel_length[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(channel_length[100]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(channel_length[101]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(channel_length[102]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(channel_length[103]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(channel_length[104]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(channel_length[105]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(channel_length[106]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(channel_length[107]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(channel_length[108]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(channel_length[109]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(channel_length[10]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(channel_length[110]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(channel_length[111]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(channel_length[112]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(channel_length[113]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(channel_length[114]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(channel_length[115]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(channel_length[116]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(channel_length[117]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(channel_length[118]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(channel_length[119]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(channel_length[11]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(channel_length[120]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(channel_length[121]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(channel_length[122]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(channel_length[123]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(channel_length[124]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(channel_length[125]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(channel_length[126]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input35 (.A(channel_length[127]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(channel_length[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(channel_length[13]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(channel_length[14]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(channel_length[15]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(channel_length[16]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(channel_length[17]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(channel_length[18]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(channel_length[19]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(channel_length[1]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(channel_length[20]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input46 (.A(channel_length[21]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input47 (.A(channel_length[22]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input48 (.A(channel_length[23]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input49 (.A(channel_length[24]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input50 (.A(channel_length[25]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input51 (.A(channel_length[26]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input52 (.A(channel_length[27]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(channel_length[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(channel_length[29]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(channel_length[2]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input56 (.A(channel_length[30]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input57 (.A(channel_length[31]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(channel_length[32]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(channel_length[33]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(channel_length[34]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(channel_length[35]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(channel_length[36]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(channel_length[37]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(channel_length[38]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(channel_length[39]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(channel_length[3]),
    .X(net67));
 sky130_fd_sc_hd__buf_6 input67 (.A(channel_length[40]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input68 (.A(channel_length[41]),
    .X(net69));
 sky130_fd_sc_hd__buf_6 input69 (.A(channel_length[42]),
    .X(net70));
 sky130_fd_sc_hd__buf_6 input70 (.A(channel_length[43]),
    .X(net71));
 sky130_fd_sc_hd__buf_6 input71 (.A(channel_length[44]),
    .X(net72));
 sky130_fd_sc_hd__buf_6 input72 (.A(channel_length[45]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_8 input73 (.A(channel_length[46]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(channel_length[47]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(channel_length[48]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(channel_length[49]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(channel_length[4]),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(channel_length[50]),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input79 (.A(channel_length[51]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(channel_length[52]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(channel_length[53]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(channel_length[54]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(channel_length[55]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(channel_length[56]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(channel_length[57]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(channel_length[58]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(channel_length[59]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(channel_length[5]),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(channel_length[60]),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(channel_length[61]),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 input91 (.A(channel_length[62]),
    .X(net92));
 sky130_fd_sc_hd__buf_6 input92 (.A(channel_length[63]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(channel_length[64]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(channel_length[65]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(channel_length[66]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(channel_length[67]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(channel_length[68]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(channel_length[69]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(channel_length[6]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(channel_length[70]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(channel_length[71]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(channel_length[72]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(channel_length[73]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(channel_length[74]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(channel_length[75]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(channel_length[76]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(channel_length[77]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(channel_length[78]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(channel_length[79]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(channel_length[7]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(channel_length[80]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(channel_length[81]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(channel_length[82]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(channel_length[83]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(channel_length[84]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(channel_length[85]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(channel_length[86]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(channel_length[87]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(channel_length[88]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(channel_length[89]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(channel_length[8]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(channel_length[90]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(channel_length[91]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(channel_length[92]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(channel_length[93]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(channel_length[94]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(channel_length[95]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(channel_length[96]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(channel_length[97]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(channel_length[98]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(channel_length[99]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(channel_length[9]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(channel_start[0]),
    .X(net134));
 sky130_fd_sc_hd__buf_2 input134 (.A(channel_start[1]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(channel_start[2]),
    .X(net136));
 sky130_fd_sc_hd__buf_4 input136 (.A(channel_start[3]),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(dst_wready[0]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(dst_wready[1]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(dst_wready[2]),
    .X(net140));
 sky130_fd_sc_hd__buf_4 input140 (.A(dst_wready[3]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(src_rvalid[0]),
    .X(net142));
 sky130_fd_sc_hd__buf_4 input142 (.A(src_rvalid[1]),
    .X(net143));
 sky130_fd_sc_hd__buf_4 input143 (.A(src_rvalid[2]),
    .X(net144));
 sky130_fd_sc_hd__buf_4 input144 (.A(src_rvalid[3]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net146),
    .X(channel_busy[0]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net147),
    .X(channel_busy[1]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net148),
    .X(channel_busy[2]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net149),
    .X(channel_busy[3]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net150),
    .X(channel_done[0]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net151),
    .X(channel_done[1]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net152),
    .X(channel_done[2]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net153),
    .X(channel_done[3]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net154),
    .X(channel_error[0]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net155),
    .X(channel_error[1]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net156),
    .X(channel_error[2]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net157),
    .X(channel_error[3]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net158),
    .X(debug_active_channels[0]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net159),
    .X(debug_active_channels[1]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net160),
    .X(debug_active_channels[2]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net161),
    .X(debug_active_channels[3]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net162),
    .X(debug_has_active_channels));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net163),
    .X(dst_write[0]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net164),
    .X(dst_write[1]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net165),
    .X(dst_write[2]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net166),
    .X(dst_write[3]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net167),
    .X(src_read[0]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net168),
    .X(src_read[1]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net169),
    .X(src_read[2]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net170),
    .X(src_read[3]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net171),
    .X(src_rready[0]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net172),
    .X(src_rready[1]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net173),
    .X(src_rready[2]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net174),
    .X(src_rready[3]));
 sky130_fd_sc_hd__conb_1 _2752__174 (.LO(net175));
 sky130_fd_sc_hd__conb_1 _2753__175 (.LO(net176));
 sky130_fd_sc_hd__conb_1 _2754__176 (.LO(net177));
 sky130_fd_sc_hd__conb_1 _2755__177 (.LO(net178));
 sky130_fd_sc_hd__conb_1 _2756__178 (.LO(net179));
 sky130_fd_sc_hd__conb_1 _2757__179 (.LO(net180));
 sky130_fd_sc_hd__conb_1 _2758__180 (.LO(net181));
 sky130_fd_sc_hd__conb_1 _2759__181 (.LO(net182));
 sky130_fd_sc_hd__conb_1 _2760__182 (.LO(net183));
 sky130_fd_sc_hd__conb_1 _2761__183 (.LO(net184));
 sky130_fd_sc_hd__conb_1 _2762__184 (.LO(net185));
 sky130_fd_sc_hd__conb_1 _2763__185 (.LO(net186));
 sky130_fd_sc_hd__conb_1 _2764__186 (.LO(net187));
 sky130_fd_sc_hd__conb_1 _2765__187 (.LO(net188));
 sky130_fd_sc_hd__conb_1 _2766__188 (.LO(net189));
 sky130_fd_sc_hd__conb_1 _2767__189 (.LO(net190));
 sky130_fd_sc_hd__conb_1 _2768__190 (.LO(net191));
 sky130_fd_sc_hd__conb_1 _2769__191 (.LO(net192));
 sky130_fd_sc_hd__conb_1 _2770__192 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _2771__193 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _2772__194 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _2773__195 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _2774__196 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _2775__197 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _2776__198 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _2777__199 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _2778__200 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _2779__201 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _2780__202 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _2781__203 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _2782__204 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _2783__205 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _2784__206 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _2785__207 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _2786__208 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _2787__209 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _2788__210 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _2789__211 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _2790__212 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _2791__213 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _2792__214 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _2793__215 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _2794__216 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _2795__217 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _2796__218 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _2797__219 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _2798__220 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _2799__221 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _2800__222 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _2801__223 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _2802__224 (.LO(net225));
 sky130_fd_sc_hd__conb_1 _2803__225 (.LO(net226));
 sky130_fd_sc_hd__conb_1 _2804__226 (.LO(net227));
 sky130_fd_sc_hd__conb_1 _2805__227 (.LO(net228));
 sky130_fd_sc_hd__conb_1 _2806__228 (.LO(net229));
 sky130_fd_sc_hd__conb_1 _2807__229 (.LO(net230));
 sky130_fd_sc_hd__conb_1 _2808__230 (.LO(net231));
 sky130_fd_sc_hd__conb_1 _2809__231 (.LO(net232));
 sky130_fd_sc_hd__conb_1 _2810__232 (.LO(net233));
 sky130_fd_sc_hd__conb_1 _2811__233 (.LO(net234));
 sky130_fd_sc_hd__conb_1 _2812__234 (.LO(net235));
 sky130_fd_sc_hd__conb_1 _2813__235 (.LO(net236));
 sky130_fd_sc_hd__conb_1 _2814__236 (.LO(net237));
 sky130_fd_sc_hd__conb_1 _2815__237 (.LO(net238));
 sky130_fd_sc_hd__conb_1 _2816__238 (.LO(net239));
 sky130_fd_sc_hd__conb_1 _2817__239 (.LO(net240));
 sky130_fd_sc_hd__conb_1 _2818__240 (.LO(net241));
 sky130_fd_sc_hd__conb_1 _2819__241 (.LO(net242));
 sky130_fd_sc_hd__conb_1 _2820__242 (.LO(net243));
 sky130_fd_sc_hd__conb_1 _2821__243 (.LO(net244));
 sky130_fd_sc_hd__conb_1 _2822__244 (.LO(net245));
 sky130_fd_sc_hd__conb_1 _2823__245 (.LO(net246));
 sky130_fd_sc_hd__conb_1 _2824__246 (.LO(net247));
 sky130_fd_sc_hd__conb_1 _2825__247 (.LO(net248));
 sky130_fd_sc_hd__conb_1 _2826__248 (.LO(net249));
 sky130_fd_sc_hd__conb_1 _2827__249 (.LO(net250));
 sky130_fd_sc_hd__conb_1 _2828__250 (.LO(net251));
 sky130_fd_sc_hd__conb_1 _2829__251 (.LO(net252));
 sky130_fd_sc_hd__conb_1 _2830__252 (.LO(net253));
 sky130_fd_sc_hd__conb_1 _2831__253 (.LO(net254));
 sky130_fd_sc_hd__conb_1 _2832__254 (.LO(net255));
 sky130_fd_sc_hd__conb_1 _2833__255 (.LO(net256));
 sky130_fd_sc_hd__conb_1 _2834__256 (.LO(net257));
 sky130_fd_sc_hd__conb_1 _2835__257 (.LO(net258));
 sky130_fd_sc_hd__conb_1 _2836__258 (.LO(net259));
 sky130_fd_sc_hd__conb_1 _2837__259 (.LO(net260));
 sky130_fd_sc_hd__conb_1 _2838__260 (.LO(net261));
 sky130_fd_sc_hd__conb_1 _2839__261 (.LO(net262));
 sky130_fd_sc_hd__conb_1 _2840__262 (.LO(net263));
 sky130_fd_sc_hd__conb_1 _2841__263 (.LO(net264));
 sky130_fd_sc_hd__conb_1 _2842__264 (.LO(net265));
 sky130_fd_sc_hd__conb_1 _2843__265 (.LO(net266));
 sky130_fd_sc_hd__conb_1 _2844__266 (.LO(net267));
 sky130_fd_sc_hd__conb_1 _2845__267 (.LO(net268));
 sky130_fd_sc_hd__conb_1 _2846__268 (.LO(net269));
 sky130_fd_sc_hd__conb_1 _2847__269 (.LO(net270));
 sky130_fd_sc_hd__conb_1 _2848__270 (.LO(net271));
 sky130_fd_sc_hd__conb_1 _2849__271 (.LO(net272));
 sky130_fd_sc_hd__conb_1 _2850__272 (.LO(net273));
 sky130_fd_sc_hd__conb_1 _2851__273 (.LO(net274));
 sky130_fd_sc_hd__conb_1 _2852__274 (.LO(net275));
 sky130_fd_sc_hd__conb_1 _2853__275 (.LO(net276));
 sky130_fd_sc_hd__conb_1 _2854__276 (.LO(net277));
 sky130_fd_sc_hd__conb_1 _2855__277 (.LO(net278));
 sky130_fd_sc_hd__conb_1 _2856__278 (.LO(net279));
 sky130_fd_sc_hd__conb_1 _2857__279 (.LO(net280));
 sky130_fd_sc_hd__conb_1 _2858__280 (.LO(net281));
 sky130_fd_sc_hd__conb_1 _2859__281 (.LO(net282));
 sky130_fd_sc_hd__conb_1 _2860__282 (.LO(net283));
 sky130_fd_sc_hd__conb_1 _2861__283 (.LO(net284));
 sky130_fd_sc_hd__conb_1 _2862__284 (.LO(net285));
 sky130_fd_sc_hd__conb_1 _2863__285 (.LO(net286));
 sky130_fd_sc_hd__conb_1 _2864__286 (.LO(net287));
 sky130_fd_sc_hd__conb_1 _2865__287 (.LO(net288));
 sky130_fd_sc_hd__conb_1 _2866__288 (.LO(net289));
 sky130_fd_sc_hd__conb_1 _2867__289 (.LO(net290));
 sky130_fd_sc_hd__conb_1 _2868__290 (.LO(net291));
 sky130_fd_sc_hd__conb_1 _2869__291 (.LO(net292));
 sky130_fd_sc_hd__conb_1 _2870__292 (.LO(net293));
 sky130_fd_sc_hd__conb_1 _2871__293 (.LO(net294));
 sky130_fd_sc_hd__conb_1 _2872__294 (.LO(net295));
 sky130_fd_sc_hd__conb_1 _2873__295 (.LO(net296));
 sky130_fd_sc_hd__conb_1 _2874__296 (.LO(net297));
 sky130_fd_sc_hd__conb_1 _2875__297 (.LO(net298));
 sky130_fd_sc_hd__conb_1 _2876__298 (.LO(net299));
 sky130_fd_sc_hd__conb_1 _2877__299 (.LO(net300));
 sky130_fd_sc_hd__conb_1 _2878__300 (.LO(net301));
 sky130_fd_sc_hd__conb_1 _2879__301 (.LO(net302));
 sky130_fd_sc_hd__conb_1 _2880__302 (.LO(net303));
 sky130_fd_sc_hd__conb_1 _2881__303 (.LO(net304));
 sky130_fd_sc_hd__conb_1 _2882__304 (.LO(net305));
 sky130_fd_sc_hd__conb_1 _2883__305 (.LO(net306));
 sky130_fd_sc_hd__conb_1 _2884__306 (.LO(net307));
 sky130_fd_sc_hd__conb_1 _2885__307 (.LO(net308));
 sky130_fd_sc_hd__conb_1 _2886__308 (.LO(net309));
 sky130_fd_sc_hd__conb_1 _2887__309 (.LO(net310));
 sky130_fd_sc_hd__conb_1 _2888__310 (.LO(net311));
 sky130_fd_sc_hd__conb_1 _2889__311 (.LO(net312));
 sky130_fd_sc_hd__conb_1 _2890__312 (.LO(net313));
 sky130_fd_sc_hd__conb_1 _2891__313 (.LO(net314));
 sky130_fd_sc_hd__conb_1 _2892__314 (.LO(net315));
 sky130_fd_sc_hd__conb_1 _2893__315 (.LO(net316));
 sky130_fd_sc_hd__conb_1 _2894__316 (.LO(net317));
 sky130_fd_sc_hd__conb_1 _2895__317 (.LO(net318));
 sky130_fd_sc_hd__conb_1 _2896__318 (.LO(net319));
 sky130_fd_sc_hd__conb_1 _2897__319 (.LO(net320));
 sky130_fd_sc_hd__conb_1 _2898__320 (.LO(net321));
 sky130_fd_sc_hd__conb_1 _2899__321 (.LO(net322));
 sky130_fd_sc_hd__conb_1 _2900__322 (.LO(net323));
 sky130_fd_sc_hd__conb_1 _2901__323 (.LO(net324));
 sky130_fd_sc_hd__conb_1 _2902__324 (.LO(net325));
 sky130_fd_sc_hd__conb_1 _2903__325 (.LO(net326));
 sky130_fd_sc_hd__conb_1 _2904__326 (.LO(net327));
 sky130_fd_sc_hd__conb_1 _2905__327 (.LO(net328));
 sky130_fd_sc_hd__conb_1 _2906__328 (.LO(net329));
 sky130_fd_sc_hd__conb_1 _2907__329 (.LO(net330));
 sky130_fd_sc_hd__conb_1 _2908__330 (.LO(net331));
 sky130_fd_sc_hd__conb_1 _2909__331 (.LO(net332));
 sky130_fd_sc_hd__conb_1 _2910__332 (.LO(net333));
 sky130_fd_sc_hd__conb_1 _2911__333 (.LO(net334));
 sky130_fd_sc_hd__conb_1 _2912__334 (.LO(net335));
 sky130_fd_sc_hd__conb_1 _2913__335 (.LO(net336));
 sky130_fd_sc_hd__conb_1 _2914__336 (.LO(net337));
 sky130_fd_sc_hd__conb_1 _2915__337 (.LO(net338));
 sky130_fd_sc_hd__conb_1 _2916__338 (.LO(net339));
 sky130_fd_sc_hd__conb_1 _2917__339 (.LO(net340));
 sky130_fd_sc_hd__conb_1 _2918__340 (.LO(net341));
 sky130_fd_sc_hd__conb_1 _2919__341 (.LO(net342));
 sky130_fd_sc_hd__conb_1 _2920__342 (.LO(net343));
 sky130_fd_sc_hd__conb_1 _2921__343 (.LO(net344));
 sky130_fd_sc_hd__conb_1 _2922__344 (.LO(net345));
 sky130_fd_sc_hd__conb_1 _2923__345 (.LO(net346));
 sky130_fd_sc_hd__conb_1 _2924__346 (.LO(net347));
 sky130_fd_sc_hd__conb_1 _2925__347 (.LO(net348));
 sky130_fd_sc_hd__conb_1 _2926__348 (.LO(net349));
 sky130_fd_sc_hd__conb_1 _2927__349 (.LO(net350));
 sky130_fd_sc_hd__conb_1 _2928__350 (.LO(net351));
 sky130_fd_sc_hd__conb_1 _2929__351 (.LO(net352));
 sky130_fd_sc_hd__conb_1 _2930__352 (.LO(net353));
 sky130_fd_sc_hd__conb_1 _2931__353 (.LO(net354));
 sky130_fd_sc_hd__conb_1 _2932__354 (.LO(net355));
 sky130_fd_sc_hd__conb_1 _2933__355 (.LO(net356));
 sky130_fd_sc_hd__conb_1 _2934__356 (.LO(net357));
 sky130_fd_sc_hd__conb_1 _2935__357 (.LO(net358));
 sky130_fd_sc_hd__conb_1 _2936__358 (.LO(net359));
 sky130_fd_sc_hd__conb_1 _2937__359 (.LO(net360));
 sky130_fd_sc_hd__conb_1 _2938__360 (.LO(net361));
 sky130_fd_sc_hd__conb_1 _2939__361 (.LO(net362));
 sky130_fd_sc_hd__conb_1 _2940__362 (.LO(net363));
 sky130_fd_sc_hd__conb_1 _2941__363 (.LO(net364));
 sky130_fd_sc_hd__conb_1 _2942__364 (.LO(net365));
 sky130_fd_sc_hd__conb_1 _2943__365 (.LO(net366));
 sky130_fd_sc_hd__conb_1 _2944__366 (.LO(net367));
 sky130_fd_sc_hd__conb_1 _2945__367 (.LO(net368));
 sky130_fd_sc_hd__conb_1 _2946__368 (.LO(net369));
 sky130_fd_sc_hd__conb_1 _2947__369 (.LO(net370));
 sky130_fd_sc_hd__conb_1 _2948__370 (.LO(net371));
 sky130_fd_sc_hd__conb_1 _2949__371 (.LO(net372));
 sky130_fd_sc_hd__conb_1 _2950__372 (.LO(net373));
 sky130_fd_sc_hd__conb_1 _2951__373 (.LO(net374));
 sky130_fd_sc_hd__conb_1 _2952__374 (.LO(net375));
 sky130_fd_sc_hd__conb_1 _2953__375 (.LO(net376));
 sky130_fd_sc_hd__conb_1 _2954__376 (.LO(net377));
 sky130_fd_sc_hd__conb_1 _2955__377 (.LO(net378));
 sky130_fd_sc_hd__conb_1 _2956__378 (.LO(net379));
 sky130_fd_sc_hd__conb_1 _2957__379 (.LO(net380));
 sky130_fd_sc_hd__conb_1 _2958__380 (.LO(net381));
 sky130_fd_sc_hd__conb_1 _2959__381 (.LO(net382));
 sky130_fd_sc_hd__conb_1 _2960__382 (.LO(net383));
 sky130_fd_sc_hd__conb_1 _2961__383 (.LO(net384));
 sky130_fd_sc_hd__conb_1 _2962__384 (.LO(net385));
 sky130_fd_sc_hd__conb_1 _2963__385 (.LO(net386));
 sky130_fd_sc_hd__conb_1 _2964__386 (.LO(net387));
 sky130_fd_sc_hd__conb_1 _2965__387 (.LO(net388));
 sky130_fd_sc_hd__conb_1 _2966__388 (.LO(net389));
 sky130_fd_sc_hd__conb_1 _2967__389 (.LO(net390));
 sky130_fd_sc_hd__conb_1 _2968__390 (.LO(net391));
 sky130_fd_sc_hd__conb_1 _2969__391 (.LO(net392));
 sky130_fd_sc_hd__conb_1 _2970__392 (.LO(net393));
 sky130_fd_sc_hd__conb_1 _2971__393 (.LO(net394));
 sky130_fd_sc_hd__conb_1 _2972__394 (.LO(net395));
 sky130_fd_sc_hd__conb_1 _2973__395 (.LO(net396));
 sky130_fd_sc_hd__conb_1 _2974__396 (.LO(net397));
 sky130_fd_sc_hd__conb_1 _2975__397 (.LO(net398));
 sky130_fd_sc_hd__conb_1 _2976__398 (.LO(net399));
 sky130_fd_sc_hd__conb_1 _2977__399 (.LO(net400));
 sky130_fd_sc_hd__conb_1 _2978__400 (.LO(net401));
 sky130_fd_sc_hd__conb_1 _2979__401 (.LO(net402));
 sky130_fd_sc_hd__conb_1 _2980__402 (.LO(net403));
 sky130_fd_sc_hd__conb_1 _2981__403 (.LO(net404));
 sky130_fd_sc_hd__conb_1 _2982__404 (.LO(net405));
 sky130_fd_sc_hd__conb_1 _2983__405 (.LO(net406));
 sky130_fd_sc_hd__conb_1 _2984__406 (.LO(net407));
 sky130_fd_sc_hd__conb_1 _2985__407 (.LO(net408));
 sky130_fd_sc_hd__conb_1 _2986__408 (.LO(net409));
 sky130_fd_sc_hd__conb_1 _2987__409 (.LO(net410));
 sky130_fd_sc_hd__conb_1 _2988__410 (.LO(net411));
 sky130_fd_sc_hd__conb_1 _2989__411 (.LO(net412));
 sky130_fd_sc_hd__conb_1 _2990__412 (.LO(net413));
 sky130_fd_sc_hd__conb_1 _2991__413 (.LO(net414));
 sky130_fd_sc_hd__conb_1 _2992__414 (.LO(net415));
 sky130_fd_sc_hd__conb_1 _2993__415 (.LO(net416));
 sky130_fd_sc_hd__conb_1 _2994__416 (.LO(net417));
 sky130_fd_sc_hd__conb_1 _2995__417 (.LO(net418));
 sky130_fd_sc_hd__conb_1 _2996__418 (.LO(net419));
 sky130_fd_sc_hd__conb_1 _2997__419 (.LO(net420));
 sky130_fd_sc_hd__conb_1 _2998__420 (.LO(net421));
 sky130_fd_sc_hd__conb_1 _2999__421 (.LO(net422));
 sky130_fd_sc_hd__conb_1 _3000__422 (.LO(net423));
 sky130_fd_sc_hd__conb_1 _3001__423 (.LO(net424));
 sky130_fd_sc_hd__conb_1 _3002__424 (.LO(net425));
 sky130_fd_sc_hd__conb_1 _3003__425 (.LO(net426));
 sky130_fd_sc_hd__conb_1 _3004__426 (.LO(net427));
 sky130_fd_sc_hd__conb_1 _3005__427 (.LO(net428));
 sky130_fd_sc_hd__conb_1 _3006__428 (.LO(net429));
 sky130_fd_sc_hd__conb_1 _3007__429 (.LO(net430));
 sky130_fd_sc_hd__conb_1 _3008__430 (.LO(net431));
 sky130_fd_sc_hd__conb_1 _3009__431 (.LO(net432));
 sky130_fd_sc_hd__conb_1 _3010__432 (.LO(net433));
 sky130_fd_sc_hd__conb_1 _3011__433 (.LO(net434));
 sky130_fd_sc_hd__conb_1 _3012__434 (.LO(net435));
 sky130_fd_sc_hd__conb_1 _3013__435 (.LO(net436));
 sky130_fd_sc_hd__conb_1 _3014__436 (.LO(net437));
 sky130_fd_sc_hd__conb_1 _3015__437 (.LO(net438));
 sky130_fd_sc_hd__conb_1 _3016__438 (.LO(net439));
 sky130_fd_sc_hd__conb_1 _3017__439 (.LO(net440));
 sky130_fd_sc_hd__conb_1 _3018__440 (.LO(net441));
 sky130_fd_sc_hd__conb_1 _3019__441 (.LO(net442));
 sky130_fd_sc_hd__conb_1 _3020__442 (.LO(net443));
 sky130_fd_sc_hd__conb_1 _3021__443 (.LO(net444));
 sky130_fd_sc_hd__conb_1 _3022__444 (.LO(net445));
 sky130_fd_sc_hd__conb_1 _3023__445 (.LO(net446));
 sky130_fd_sc_hd__conb_1 _3024__446 (.LO(net447));
 sky130_fd_sc_hd__conb_1 _3025__447 (.LO(net448));
 sky130_fd_sc_hd__conb_1 _3026__448 (.LO(net449));
 sky130_fd_sc_hd__conb_1 _3027__449 (.LO(net450));
 sky130_fd_sc_hd__conb_1 _3028__450 (.LO(net451));
 sky130_fd_sc_hd__conb_1 _3029__451 (.LO(net452));
 sky130_fd_sc_hd__conb_1 _3030__452 (.LO(net453));
 sky130_fd_sc_hd__conb_1 _3031__453 (.LO(net454));
 sky130_fd_sc_hd__conb_1 _3032__454 (.LO(net455));
 sky130_fd_sc_hd__conb_1 _3033__455 (.LO(net456));
 sky130_fd_sc_hd__conb_1 _3034__456 (.LO(net457));
 sky130_fd_sc_hd__conb_1 _3035__457 (.LO(net458));
 sky130_fd_sc_hd__conb_1 _3036__458 (.LO(net459));
 sky130_fd_sc_hd__conb_1 _3037__459 (.LO(net460));
 sky130_fd_sc_hd__conb_1 _3038__460 (.LO(net461));
 sky130_fd_sc_hd__conb_1 _3039__461 (.LO(net462));
 sky130_fd_sc_hd__conb_1 _3040__462 (.LO(net463));
 sky130_fd_sc_hd__conb_1 _3041__463 (.LO(net464));
 sky130_fd_sc_hd__conb_1 _3042__464 (.LO(net465));
 sky130_fd_sc_hd__conb_1 _3043__465 (.LO(net466));
 sky130_fd_sc_hd__conb_1 _3044__466 (.LO(net467));
 sky130_fd_sc_hd__conb_1 _3045__467 (.LO(net468));
 sky130_fd_sc_hd__conb_1 _3046__468 (.LO(net469));
 sky130_fd_sc_hd__conb_1 _3047__469 (.LO(net470));
 sky130_fd_sc_hd__conb_1 _3048__470 (.LO(net471));
 sky130_fd_sc_hd__conb_1 _3049__471 (.LO(net472));
 sky130_fd_sc_hd__conb_1 _3050__472 (.LO(net473));
 sky130_fd_sc_hd__conb_1 _3051__473 (.LO(net474));
 sky130_fd_sc_hd__conb_1 _3052__474 (.LO(net475));
 sky130_fd_sc_hd__conb_1 _3053__475 (.LO(net476));
 sky130_fd_sc_hd__conb_1 _3054__476 (.LO(net477));
 sky130_fd_sc_hd__conb_1 _3055__477 (.LO(net478));
 sky130_fd_sc_hd__conb_1 _3056__478 (.LO(net479));
 sky130_fd_sc_hd__conb_1 _3057__479 (.LO(net480));
 sky130_fd_sc_hd__conb_1 _3058__480 (.LO(net481));
 sky130_fd_sc_hd__conb_1 _3059__481 (.LO(net482));
 sky130_fd_sc_hd__conb_1 _3060__482 (.LO(net483));
 sky130_fd_sc_hd__conb_1 _3061__483 (.LO(net484));
 sky130_fd_sc_hd__conb_1 _3062__484 (.LO(net485));
 sky130_fd_sc_hd__conb_1 _3063__485 (.LO(net486));
 sky130_fd_sc_hd__conb_1 _3064__486 (.LO(net487));
 sky130_fd_sc_hd__conb_1 _3065__487 (.LO(net488));
 sky130_fd_sc_hd__conb_1 _3066__488 (.LO(net489));
 sky130_fd_sc_hd__conb_1 _3067__489 (.LO(net490));
 sky130_fd_sc_hd__conb_1 _3068__490 (.LO(net491));
 sky130_fd_sc_hd__conb_1 _3069__491 (.LO(net492));
 sky130_fd_sc_hd__conb_1 _3070__492 (.LO(net493));
 sky130_fd_sc_hd__conb_1 _3071__493 (.LO(net494));
 sky130_fd_sc_hd__conb_1 _3072__494 (.LO(net495));
 sky130_fd_sc_hd__conb_1 _3073__495 (.LO(net496));
 sky130_fd_sc_hd__conb_1 _3074__496 (.LO(net497));
 sky130_fd_sc_hd__conb_1 _3075__497 (.LO(net498));
 sky130_fd_sc_hd__conb_1 _3076__498 (.LO(net499));
 sky130_fd_sc_hd__conb_1 _3077__499 (.LO(net500));
 sky130_fd_sc_hd__conb_1 _3078__500 (.LO(net501));
 sky130_fd_sc_hd__conb_1 _3079__501 (.LO(net502));
 sky130_fd_sc_hd__conb_1 _3080__502 (.LO(net503));
 sky130_fd_sc_hd__conb_1 _3081__503 (.LO(net504));
 sky130_fd_sc_hd__conb_1 _3082__504 (.LO(net505));
 sky130_fd_sc_hd__conb_1 _3083__505 (.LO(net506));
 sky130_fd_sc_hd__conb_1 _3084__506 (.LO(net507));
 sky130_fd_sc_hd__conb_1 _3085__507 (.LO(net508));
 sky130_fd_sc_hd__conb_1 _3086__508 (.LO(net509));
 sky130_fd_sc_hd__conb_1 _3087__509 (.LO(net510));
 sky130_fd_sc_hd__conb_1 _3088__510 (.LO(net511));
 sky130_fd_sc_hd__conb_1 _3089__511 (.LO(net512));
 sky130_fd_sc_hd__conb_1 _3090__512 (.LO(net513));
 sky130_fd_sc_hd__conb_1 _3091__513 (.LO(net514));
 sky130_fd_sc_hd__conb_1 _3092__514 (.LO(net515));
 sky130_fd_sc_hd__conb_1 _3093__515 (.LO(net516));
 sky130_fd_sc_hd__conb_1 _3094__516 (.LO(net517));
 sky130_fd_sc_hd__conb_1 _3095__517 (.LO(net518));
 sky130_fd_sc_hd__conb_1 _3096__518 (.LO(net519));
 sky130_fd_sc_hd__conb_1 _3097__519 (.LO(net520));
 sky130_fd_sc_hd__conb_1 _3098__520 (.LO(net521));
 sky130_fd_sc_hd__conb_1 _3099__521 (.LO(net522));
 sky130_fd_sc_hd__conb_1 _3100__522 (.LO(net523));
 sky130_fd_sc_hd__conb_1 _3101__523 (.LO(net524));
 sky130_fd_sc_hd__conb_1 _3102__524 (.LO(net525));
 sky130_fd_sc_hd__conb_1 _3103__525 (.LO(net526));
 sky130_fd_sc_hd__conb_1 _3104__526 (.LO(net527));
 sky130_fd_sc_hd__conb_1 _3105__527 (.LO(net528));
 sky130_fd_sc_hd__conb_1 _3106__528 (.LO(net529));
 sky130_fd_sc_hd__conb_1 _3107__529 (.LO(net530));
 sky130_fd_sc_hd__conb_1 _3108__530 (.LO(net531));
 sky130_fd_sc_hd__conb_1 _3109__531 (.LO(net532));
 sky130_fd_sc_hd__conb_1 _3110__532 (.LO(net533));
 sky130_fd_sc_hd__conb_1 _3111__533 (.LO(net534));
 sky130_fd_sc_hd__conb_1 _3112__534 (.LO(net535));
 sky130_fd_sc_hd__conb_1 _3113__535 (.LO(net536));
 sky130_fd_sc_hd__conb_1 _3114__536 (.LO(net537));
 sky130_fd_sc_hd__conb_1 _3115__537 (.LO(net538));
 sky130_fd_sc_hd__conb_1 _3116__538 (.LO(net539));
 sky130_fd_sc_hd__conb_1 _3117__539 (.LO(net540));
 sky130_fd_sc_hd__conb_1 _3118__540 (.LO(net541));
 sky130_fd_sc_hd__conb_1 _3119__541 (.LO(net542));
 sky130_fd_sc_hd__conb_1 _3120__542 (.LO(net543));
 sky130_fd_sc_hd__conb_1 _3121__543 (.LO(net544));
 sky130_fd_sc_hd__conb_1 _3122__544 (.LO(net545));
 sky130_fd_sc_hd__conb_1 _3123__545 (.LO(net546));
 sky130_fd_sc_hd__conb_1 _3124__546 (.LO(net547));
 sky130_fd_sc_hd__conb_1 _3125__547 (.LO(net548));
 sky130_fd_sc_hd__conb_1 _3126__548 (.LO(net549));
 sky130_fd_sc_hd__conb_1 _3127__549 (.LO(net550));
 sky130_fd_sc_hd__conb_1 _3128__550 (.LO(net551));
 sky130_fd_sc_hd__conb_1 _3129__551 (.LO(net552));
 sky130_fd_sc_hd__conb_1 _3130__552 (.LO(net553));
 sky130_fd_sc_hd__conb_1 _3131__553 (.LO(net554));
 sky130_fd_sc_hd__conb_1 _3132__554 (.LO(net555));
 sky130_fd_sc_hd__conb_1 _3133__555 (.LO(net556));
 sky130_fd_sc_hd__conb_1 _3134__556 (.LO(net557));
 sky130_fd_sc_hd__conb_1 _3135__557 (.LO(net558));
 sky130_fd_sc_hd__conb_1 _3136__558 (.LO(net559));
 sky130_fd_sc_hd__conb_1 _3137__559 (.LO(net560));
 sky130_fd_sc_hd__conb_1 _3138__560 (.LO(net561));
 sky130_fd_sc_hd__conb_1 _3139__561 (.LO(net562));
 sky130_fd_sc_hd__conb_1 _3140__562 (.LO(net563));
 sky130_fd_sc_hd__conb_1 _3141__563 (.LO(net564));
 sky130_fd_sc_hd__conb_1 _3142__564 (.LO(net565));
 sky130_fd_sc_hd__conb_1 _3143__565 (.LO(net566));
 sky130_fd_sc_hd__conb_1 _3144__566 (.LO(net567));
 sky130_fd_sc_hd__conb_1 _3145__567 (.LO(net568));
 sky130_fd_sc_hd__conb_1 _3146__568 (.LO(net569));
 sky130_fd_sc_hd__conb_1 _3147__569 (.LO(net570));
 sky130_fd_sc_hd__conb_1 _3148__570 (.LO(net571));
 sky130_fd_sc_hd__conb_1 _3149__571 (.LO(net572));
 sky130_fd_sc_hd__conb_1 _3150__572 (.LO(net573));
 sky130_fd_sc_hd__conb_1 _3151__573 (.LO(net574));
 sky130_fd_sc_hd__conb_1 _3152__574 (.LO(net575));
 sky130_fd_sc_hd__conb_1 _3153__575 (.LO(net576));
 sky130_fd_sc_hd__conb_1 _3154__576 (.LO(net577));
 sky130_fd_sc_hd__conb_1 _3155__577 (.LO(net578));
 sky130_fd_sc_hd__conb_1 _3156__578 (.LO(net579));
 sky130_fd_sc_hd__conb_1 _3157__579 (.LO(net580));
 sky130_fd_sc_hd__conb_1 _3158__580 (.LO(net581));
 sky130_fd_sc_hd__conb_1 _3159__581 (.LO(net582));
 sky130_fd_sc_hd__conb_1 _3160__582 (.LO(net583));
 sky130_fd_sc_hd__conb_1 _3161__583 (.LO(net584));
 sky130_fd_sc_hd__conb_1 _3162__584 (.LO(net585));
 sky130_fd_sc_hd__conb_1 _3163__585 (.LO(net586));
 sky130_fd_sc_hd__conb_1 _3164__586 (.LO(net587));
 sky130_fd_sc_hd__conb_1 _3165__587 (.LO(net588));
 sky130_fd_sc_hd__conb_1 _3166__588 (.LO(net589));
 sky130_fd_sc_hd__conb_1 _3167__589 (.LO(net590));
 sky130_fd_sc_hd__conb_1 _3168__590 (.LO(net591));
 sky130_fd_sc_hd__conb_1 _3169__591 (.LO(net592));
 sky130_fd_sc_hd__conb_1 _3170__592 (.LO(net593));
 sky130_fd_sc_hd__conb_1 _3171__593 (.LO(net594));
 sky130_fd_sc_hd__conb_1 _3172__594 (.LO(net595));
 sky130_fd_sc_hd__conb_1 _3173__595 (.LO(net596));
 sky130_fd_sc_hd__conb_1 _3174__596 (.LO(net597));
 sky130_fd_sc_hd__conb_1 _3175__597 (.LO(net598));
 sky130_fd_sc_hd__conb_1 _3176__598 (.LO(net599));
 sky130_fd_sc_hd__conb_1 _3177__599 (.LO(net600));
 sky130_fd_sc_hd__conb_1 _3178__600 (.LO(net601));
 sky130_fd_sc_hd__conb_1 _3179__601 (.LO(net602));
 sky130_fd_sc_hd__conb_1 _3180__602 (.LO(net603));
 sky130_fd_sc_hd__conb_1 _3181__603 (.LO(net604));
 sky130_fd_sc_hd__conb_1 _3182__604 (.LO(net605));
 sky130_fd_sc_hd__conb_1 _3183__605 (.LO(net606));
 sky130_fd_sc_hd__conb_1 _3184__606 (.LO(net607));
 sky130_fd_sc_hd__conb_1 _3185__607 (.LO(net608));
 sky130_fd_sc_hd__conb_1 _3186__608 (.LO(net609));
 sky130_fd_sc_hd__conb_1 _3187__609 (.LO(net610));
 sky130_fd_sc_hd__conb_1 _3188__610 (.LO(net611));
 sky130_fd_sc_hd__conb_1 _3189__611 (.LO(net612));
 sky130_fd_sc_hd__conb_1 _3190__612 (.LO(net613));
 sky130_fd_sc_hd__conb_1 _3191__613 (.LO(net614));
 sky130_fd_sc_hd__conb_1 _3192__614 (.LO(net615));
 sky130_fd_sc_hd__conb_1 _3193__615 (.LO(net616));
 sky130_fd_sc_hd__conb_1 _3194__616 (.LO(net617));
 sky130_fd_sc_hd__conb_1 _3195__617 (.LO(net618));
 sky130_fd_sc_hd__conb_1 _3196__618 (.LO(net619));
 sky130_fd_sc_hd__conb_1 _3197__619 (.LO(net620));
 sky130_fd_sc_hd__conb_1 _3198__620 (.LO(net621));
 sky130_fd_sc_hd__conb_1 _3199__621 (.LO(net622));
 sky130_fd_sc_hd__conb_1 _3200__622 (.LO(net623));
 sky130_fd_sc_hd__conb_1 _3201__623 (.LO(net624));
 sky130_fd_sc_hd__conb_1 _3202__624 (.LO(net625));
 sky130_fd_sc_hd__conb_1 _3203__625 (.LO(net626));
 sky130_fd_sc_hd__conb_1 _3204__626 (.LO(net627));
 sky130_fd_sc_hd__conb_1 _3205__627 (.LO(net628));
 sky130_fd_sc_hd__conb_1 _3206__628 (.LO(net629));
 sky130_fd_sc_hd__conb_1 _3207__629 (.LO(net630));
 sky130_fd_sc_hd__conb_1 _3208__630 (.LO(net631));
 sky130_fd_sc_hd__conb_1 _3209__631 (.LO(net632));
 sky130_fd_sc_hd__conb_1 _3210__632 (.LO(net633));
 sky130_fd_sc_hd__conb_1 _3211__633 (.LO(net634));
 sky130_fd_sc_hd__conb_1 _3212__634 (.LO(net635));
 sky130_fd_sc_hd__conb_1 _3213__635 (.LO(net636));
 sky130_fd_sc_hd__conb_1 _3214__636 (.LO(net637));
 sky130_fd_sc_hd__conb_1 _3215__637 (.LO(net638));
 sky130_fd_sc_hd__conb_1 _3216__638 (.LO(net639));
 sky130_fd_sc_hd__conb_1 _3217__639 (.LO(net640));
 sky130_fd_sc_hd__conb_1 _3218__640 (.LO(net641));
 sky130_fd_sc_hd__conb_1 _3219__641 (.LO(net642));
 sky130_fd_sc_hd__conb_1 _3220__642 (.LO(net643));
 sky130_fd_sc_hd__conb_1 _3221__643 (.LO(net644));
 sky130_fd_sc_hd__conb_1 _3222__644 (.LO(net645));
 sky130_fd_sc_hd__conb_1 _3223__645 (.LO(net646));
 sky130_fd_sc_hd__conb_1 _3224__646 (.LO(net647));
 sky130_fd_sc_hd__conb_1 _3225__647 (.LO(net648));
 sky130_fd_sc_hd__conb_1 _3226__648 (.LO(net649));
 sky130_fd_sc_hd__conb_1 _3227__649 (.LO(net650));
 sky130_fd_sc_hd__conb_1 _3228__650 (.LO(net651));
 sky130_fd_sc_hd__conb_1 _3229__651 (.LO(net652));
 sky130_fd_sc_hd__conb_1 _3230__652 (.LO(net653));
 sky130_fd_sc_hd__conb_1 _3231__653 (.LO(net654));
 sky130_fd_sc_hd__conb_1 _3232__654 (.LO(net655));
 sky130_fd_sc_hd__conb_1 _3233__655 (.LO(net656));
 sky130_fd_sc_hd__conb_1 _3234__656 (.LO(net657));
 sky130_fd_sc_hd__conb_1 _3235__657 (.LO(net658));
 sky130_fd_sc_hd__conb_1 _3236__658 (.LO(net659));
 sky130_fd_sc_hd__conb_1 _3237__659 (.LO(net660));
 sky130_fd_sc_hd__conb_1 _3238__660 (.LO(net661));
 sky130_fd_sc_hd__conb_1 _3239__661 (.LO(net662));
 sky130_fd_sc_hd__conb_1 _3240__662 (.LO(net663));
 sky130_fd_sc_hd__conb_1 _3241__663 (.LO(net664));
 sky130_fd_sc_hd__conb_1 _3242__664 (.LO(net665));
 sky130_fd_sc_hd__conb_1 _3243__665 (.LO(net666));
 sky130_fd_sc_hd__conb_1 _3244__666 (.LO(net667));
 sky130_fd_sc_hd__conb_1 _3245__667 (.LO(net668));
 sky130_fd_sc_hd__conb_1 _3246__668 (.LO(net669));
 sky130_fd_sc_hd__conb_1 _3247__669 (.LO(net670));
 sky130_fd_sc_hd__conb_1 _3248__670 (.LO(net671));
 sky130_fd_sc_hd__conb_1 _3249__671 (.LO(net672));
 sky130_fd_sc_hd__conb_1 _3250__672 (.LO(net673));
 sky130_fd_sc_hd__conb_1 _3251__673 (.LO(net674));
 sky130_fd_sc_hd__conb_1 _3252__674 (.LO(net675));
 sky130_fd_sc_hd__conb_1 _3253__675 (.LO(net676));
 sky130_fd_sc_hd__conb_1 _3254__676 (.LO(net677));
 sky130_fd_sc_hd__conb_1 _3255__677 (.LO(net678));
 sky130_fd_sc_hd__conb_1 _3256__678 (.LO(net679));
 sky130_fd_sc_hd__conb_1 _3257__679 (.LO(net680));
 sky130_fd_sc_hd__conb_1 _3258__680 (.LO(net681));
 sky130_fd_sc_hd__conb_1 _3259__681 (.LO(net682));
 sky130_fd_sc_hd__conb_1 _3260__682 (.LO(net683));
 sky130_fd_sc_hd__conb_1 _3261__683 (.LO(net684));
 sky130_fd_sc_hd__conb_1 _3262__684 (.LO(net685));
 sky130_fd_sc_hd__conb_1 _3263__685 (.LO(net686));
 sky130_fd_sc_hd__conb_1 _3264__686 (.LO(net687));
 sky130_fd_sc_hd__conb_1 _3265__687 (.LO(net688));
 sky130_fd_sc_hd__conb_1 _3266__688 (.LO(net689));
 sky130_fd_sc_hd__conb_1 _3267__689 (.LO(net690));
 sky130_fd_sc_hd__conb_1 _3268__690 (.LO(net691));
 sky130_fd_sc_hd__conb_1 _3269__691 (.LO(net692));
 sky130_fd_sc_hd__conb_1 _3270__692 (.LO(net693));
 sky130_fd_sc_hd__conb_1 _3271__693 (.LO(net694));
 sky130_fd_sc_hd__conb_1 _3272__694 (.LO(net695));
 sky130_fd_sc_hd__conb_1 _3273__695 (.LO(net696));
 sky130_fd_sc_hd__conb_1 _3274__696 (.LO(net697));
 sky130_fd_sc_hd__conb_1 _3275__697 (.LO(net698));
 sky130_fd_sc_hd__conb_1 _3276__698 (.LO(net699));
 sky130_fd_sc_hd__conb_1 _3277__699 (.LO(net700));
 sky130_fd_sc_hd__conb_1 _3278__700 (.LO(net701));
 sky130_fd_sc_hd__conb_1 _3279__701 (.LO(net702));
 sky130_fd_sc_hd__conb_1 _3280__702 (.LO(net703));
 sky130_fd_sc_hd__conb_1 _3281__703 (.LO(net704));
 sky130_fd_sc_hd__conb_1 _3282__704 (.LO(net705));
 sky130_fd_sc_hd__conb_1 _3283__705 (.LO(net706));
 sky130_fd_sc_hd__conb_1 _3284__706 (.LO(net707));
 sky130_fd_sc_hd__conb_1 _3285__707 (.LO(net708));
 sky130_fd_sc_hd__conb_1 _3286__708 (.LO(net709));
 sky130_fd_sc_hd__conb_1 _3287__709 (.LO(net710));
 sky130_fd_sc_hd__conb_1 _3288__710 (.LO(net711));
 sky130_fd_sc_hd__conb_1 _3289__711 (.LO(net712));
 sky130_fd_sc_hd__conb_1 _3290__712 (.LO(net713));
 sky130_fd_sc_hd__conb_1 _3291__713 (.LO(net714));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_12 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_12 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_12 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_12 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_8 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_6 clkload13 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_1442_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_889 ();
endmodule
