module configurable_conditional_sum_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sky130_fd_sc_hd__inv_1 _249_ (.A(net13),
    .Y(_155_));
 sky130_fd_sc_hd__inv_1 _250_ (.A(net17),
    .Y(_161_));
 sky130_fd_sc_hd__inv_1 _251_ (.A(net21),
    .Y(_167_));
 sky130_fd_sc_hd__inv_1 _252_ (.A(net27),
    .Y(_173_));
 sky130_fd_sc_hd__inv_1 _253_ (.A(net31),
    .Y(_227_));
 sky130_fd_sc_hd__inv_1 _254_ (.A(net4),
    .Y(_233_));
 sky130_fd_sc_hd__inv_1 _255_ (.A(net1),
    .Y(_239_));
 sky130_fd_sc_hd__inv_1 _256_ (.A(net8),
    .Y(_245_));
 sky130_fd_sc_hd__inv_1 _257_ (.A(net45),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _258_ (.A(net49),
    .Y(_162_));
 sky130_fd_sc_hd__inv_1 _259_ (.A(net53),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _260_ (.A(net59),
    .Y(_174_));
 sky130_fd_sc_hd__inv_1 _261_ (.A(net63),
    .Y(_228_));
 sky130_fd_sc_hd__inv_1 _262_ (.A(net36),
    .Y(_234_));
 sky130_fd_sc_hd__inv_1 _263_ (.A(net33),
    .Y(_240_));
 sky130_fd_sc_hd__inv_1 _264_ (.A(net40),
    .Y(_246_));
 sky130_fd_sc_hd__or2_0 _265_ (.A(net22),
    .B(net54),
    .X(_000_));
 sky130_fd_sc_hd__inv_1 _266_ (.A(_207_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(net9),
    .B(net41),
    .Y(_002_));
 sky130_fd_sc_hd__or2_0 _268_ (.A(_247_),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__nor2_1 _269_ (.A(net10),
    .B(net42),
    .Y(_004_));
 sky130_fd_sc_hd__a21oi_1 _270_ (.A1(_001_),
    .A2(_003_),
    .B1(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__o22a_1 _271_ (.A1(net11),
    .A2(net43),
    .B1(_205_),
    .B2(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nor2_1 _272_ (.A(_203_),
    .B(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _273_ (.A(net14),
    .B(net46),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_1 _274_ (.A(_157_),
    .B(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__o22a_1 _275_ (.A1(net15),
    .A2(net47),
    .B1(_213_),
    .B2(_009_),
    .X(_010_));
 sky130_fd_sc_hd__nor3_1 _276_ (.A(_211_),
    .B(_007_),
    .C(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2b_1 _277_ (.A(_008_),
    .B_N(_159_),
    .Y(_012_));
 sky130_fd_sc_hd__o22a_1 _278_ (.A1(net15),
    .A2(net47),
    .B1(_213_),
    .B2(_012_),
    .X(_013_));
 sky130_fd_sc_hd__nor4_1 _279_ (.A(_203_),
    .B(_211_),
    .C(_013_),
    .D(_006_),
    .Y(_014_));
 sky130_fd_sc_hd__or2_1 _280_ (.A(net26),
    .B(net58),
    .X(_015_));
 sky130_fd_sc_hd__nand2b_1 _281_ (.A_N(_241_),
    .B(net65),
    .Y(_016_));
 sky130_fd_sc_hd__or2b_1 _282_ (.A(net65),
    .B_N(_243_),
    .X(_017_));
 sky130_fd_sc_hd__o22ai_1 _283_ (.A1(net12),
    .A2(net44),
    .B1(net23),
    .B2(net55),
    .Y(_018_));
 sky130_fd_sc_hd__a21oi_1 _284_ (.A1(_016_),
    .A2(_017_),
    .B1(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net23),
    .A2(net55),
    .B1(_183_),
    .X(_020_));
 sky130_fd_sc_hd__or3_2 _286_ (.A(_181_),
    .B(_019_),
    .C(_020_),
    .X(_021_));
 sky130_fd_sc_hd__a21oi_4 _287_ (.A1(_015_),
    .A2(_021_),
    .B1(_179_),
    .Y(_022_));
 sky130_fd_sc_hd__o21ai_0 _288_ (.A1(net29),
    .A2(net61),
    .B1(_189_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2b_1 _289_ (.A_N(_187_),
    .B(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__o22ai_2 _290_ (.A1(net28),
    .A2(net60),
    .B1(net29),
    .B2(net61),
    .Y(_025_));
 sky130_fd_sc_hd__nor2_1 _291_ (.A(_175_),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__o22a_1 _292_ (.A1(net30),
    .A2(net62),
    .B1(_179_),
    .B2(_015_),
    .X(_027_));
 sky130_fd_sc_hd__o21a_1 _293_ (.A1(_024_),
    .A2(_026_),
    .B1(_027_),
    .X(_028_));
 sky130_fd_sc_hd__or2_0 _294_ (.A(_185_),
    .B(_028_),
    .X(_029_));
 sky130_fd_sc_hd__or2_0 _295_ (.A(net3),
    .B(net35),
    .X(_030_));
 sky130_fd_sc_hd__o21ai_1 _296_ (.A1(net2),
    .A2(net34),
    .B1(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_1 _297_ (.A(_229_),
    .Y(_032_));
 sky130_fd_sc_hd__or2_0 _298_ (.A(net32),
    .B(net64),
    .X(_033_));
 sky130_fd_sc_hd__a21oi_1 _299_ (.A1(_032_),
    .A2(_033_),
    .B1(_195_),
    .Y(_034_));
 sky130_fd_sc_hd__a21oi_1 _300_ (.A1(_193_),
    .A2(_030_),
    .B1(_191_),
    .Y(_035_));
 sky130_fd_sc_hd__o21a_1 _301_ (.A1(_031_),
    .A2(_034_),
    .B1(_035_),
    .X(_036_));
 sky130_fd_sc_hd__inv_1 _302_ (.A(_201_),
    .Y(_037_));
 sky130_fd_sc_hd__o21bai_1 _303_ (.A1(net5),
    .A2(net37),
    .B1_N(_235_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _304_ (.A(net6),
    .B(net38),
    .Y(_039_));
 sky130_fd_sc_hd__a21oi_1 _305_ (.A1(_037_),
    .A2(_038_),
    .B1(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__o22a_1 _306_ (.A1(net7),
    .A2(net39),
    .B1(_199_),
    .B2(_040_),
    .X(_041_));
 sky130_fd_sc_hd__nor3_1 _307_ (.A(_197_),
    .B(_036_),
    .C(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__o21ai_0 _308_ (.A1(net5),
    .A2(net37),
    .B1(_237_),
    .Y(_043_));
 sky130_fd_sc_hd__a21oi_1 _309_ (.A1(_037_),
    .A2(_043_),
    .B1(_039_),
    .Y(_044_));
 sky130_fd_sc_hd__o22a_1 _310_ (.A1(net7),
    .A2(net39),
    .B1(_199_),
    .B2(_044_),
    .X(_045_));
 sky130_fd_sc_hd__nor3b_1 _311_ (.A(_197_),
    .B(_045_),
    .C_N(_036_),
    .Y(_046_));
 sky130_fd_sc_hd__or4_1 _312_ (.A(_179_),
    .B(_181_),
    .C(_019_),
    .D(_020_),
    .X(_047_));
 sky130_fd_sc_hd__inv_1 _313_ (.A(_177_),
    .Y(_048_));
 sky130_fd_sc_hd__nor2_1 _314_ (.A(_048_),
    .B(_025_),
    .Y(_049_));
 sky130_fd_sc_hd__o22a_1 _315_ (.A1(net30),
    .A2(net62),
    .B1(_024_),
    .B2(_049_),
    .X(_050_));
 sky130_fd_sc_hd__a211o_1 _316_ (.A1(_028_),
    .A2(_047_),
    .B1(_050_),
    .C1(_185_),
    .X(_051_));
 sky130_fd_sc_hd__o221ai_2 _317_ (.A1(_022_),
    .A2(_029_),
    .B1(_042_),
    .B2(_046_),
    .C1(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _318_ (.A1(_028_),
    .A2(_047_),
    .B1(_050_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_1 _319_ (.A(_179_),
    .Y(_054_));
 sky130_fd_sc_hd__o31ai_1 _320_ (.A1(_181_),
    .A2(_019_),
    .A3(_020_),
    .B1(_015_),
    .Y(_055_));
 sky130_fd_sc_hd__a21oi_1 _321_ (.A1(_054_),
    .A2(_055_),
    .B1(_028_),
    .Y(_056_));
 sky130_fd_sc_hd__a21oi_1 _322_ (.A1(_231_),
    .A2(_033_),
    .B1(_195_),
    .Y(_057_));
 sky130_fd_sc_hd__o21a_1 _323_ (.A1(_031_),
    .A2(_057_),
    .B1(_035_),
    .X(_058_));
 sky130_fd_sc_hd__nor3_1 _324_ (.A(_197_),
    .B(_058_),
    .C(_041_),
    .Y(_059_));
 sky130_fd_sc_hd__nor3b_1 _325_ (.A(_197_),
    .B(_045_),
    .C_N(_058_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_1 _326_ (.A(_185_),
    .Y(_061_));
 sky130_fd_sc_hd__o221ai_2 _327_ (.A1(_053_),
    .A2(_056_),
    .B1(_059_),
    .B2(_060_),
    .C1(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__and2_0 _328_ (.A(_052_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__buf_6 _329_ (.A(_063_),
    .X(_064_));
 sky130_fd_sc_hd__o21ai_1 _330_ (.A1(_011_),
    .A2(_014_),
    .B1(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__o21ai_0 _331_ (.A1(net9),
    .A2(net41),
    .B1(_153_),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_1 _332_ (.A1(_001_),
    .A2(_066_),
    .B1(_004_),
    .Y(_067_));
 sky130_fd_sc_hd__o22a_1 _333_ (.A1(net11),
    .A2(net43),
    .B1(_205_),
    .B2(_067_),
    .X(_068_));
 sky130_fd_sc_hd__nor2_1 _334_ (.A(_203_),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__or3_1 _335_ (.A(_211_),
    .B(_069_),
    .C(_010_),
    .X(_070_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(_211_),
    .B(_013_),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_1 _337_ (.A(_069_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__a21o_1 _338_ (.A1(_070_),
    .A2(_072_),
    .B1(_064_),
    .X(_073_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_065_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_1 _340_ (.A(net18),
    .B(net50),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(_163_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__o22a_1 _342_ (.A1(net19),
    .A2(net51),
    .B1(_219_),
    .B2(_076_),
    .X(_077_));
 sky130_fd_sc_hd__nor2_1 _343_ (.A(_217_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(net20),
    .B(net52),
    .Y(_079_));
 sky130_fd_sc_hd__o21ba_1 _345_ (.A1(_078_),
    .A2(_079_),
    .B1_N(_215_),
    .X(_080_));
 sky130_fd_sc_hd__and2_0 _346_ (.A(_171_),
    .B(_080_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _347_ (.A(_169_),
    .B(_080_),
    .Y(_082_));
 sky130_fd_sc_hd__or2_1 _348_ (.A(net16),
    .B(net48),
    .X(_083_));
 sky130_fd_sc_hd__o21ai_1 _349_ (.A1(_081_),
    .A2(_082_),
    .B1(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__o22ai_1 _350_ (.A1(net15),
    .A2(net47),
    .B1(_213_),
    .B2(_012_),
    .Y(_085_));
 sky130_fd_sc_hd__nand3_1 _351_ (.A(_052_),
    .B(_062_),
    .C(_007_),
    .Y(_086_));
 sky130_fd_sc_hd__o31a_1 _352_ (.A1(_203_),
    .A2(_068_),
    .A3(_064_),
    .B1(_086_),
    .X(_087_));
 sky130_fd_sc_hd__o311ai_2 _353_ (.A1(_203_),
    .A2(_068_),
    .A3(_064_),
    .B1(_086_),
    .C1(_010_),
    .Y(_088_));
 sky130_fd_sc_hd__nor2b_1 _354_ (.A(_075_),
    .B_N(_165_),
    .Y(_089_));
 sky130_fd_sc_hd__o22a_1 _355_ (.A1(net19),
    .A2(net51),
    .B1(_219_),
    .B2(_089_),
    .X(_090_));
 sky130_fd_sc_hd__nor2_1 _356_ (.A(_217_),
    .B(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__o21bai_1 _357_ (.A1(_079_),
    .A2(_091_),
    .B1_N(_215_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _358_ (.A(_171_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__a2111oi_1 _359_ (.A1(_169_),
    .A2(_092_),
    .B1(_093_),
    .C1(_209_),
    .D1(_211_),
    .Y(_094_));
 sky130_fd_sc_hd__o211ai_2 _360_ (.A1(_085_),
    .A2(_087_),
    .B1(_088_),
    .C1(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__nor2_1 _361_ (.A(_079_),
    .B(_091_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _362_ (.A(_215_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _363_ (.A(_209_),
    .B(_083_),
    .Y(_098_));
 sky130_fd_sc_hd__a22o_1 _364_ (.A1(_209_),
    .A2(_080_),
    .B1(_097_),
    .B2(_098_),
    .X(_099_));
 sky130_fd_sc_hd__nand2b_1 _365_ (.A_N(_080_),
    .B(_209_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_092_),
    .B(_098_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_1 _367_ (.A1(_100_),
    .A2(_101_),
    .B1(_169_),
    .Y(_102_));
 sky130_fd_sc_hd__a21oi_1 _368_ (.A1(_171_),
    .A2(_099_),
    .B1(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__o211ai_4 _369_ (.A1(_074_),
    .A2(_084_),
    .B1(_095_),
    .C1(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _370_ (.A1(_000_),
    .A2(_104_),
    .B1(_225_),
    .Y(_105_));
 sky130_fd_sc_hd__or2_0 _371_ (.A(net25),
    .B(net57),
    .X(_106_));
 sky130_fd_sc_hd__o21ai_0 _372_ (.A1(net24),
    .A2(net56),
    .B1(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _373_ (.A1(_223_),
    .A2(_106_),
    .B1(_221_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_0 _374_ (.A1(_105_),
    .A2(_107_),
    .B1(_108_),
    .Y(net66));
 sky130_fd_sc_hd__xor2_1 _375_ (.A(net65),
    .B(_242_),
    .X(net67));
 sky130_fd_sc_hd__o21ai_2 _376_ (.A1(_022_),
    .A2(_029_),
    .B1(_051_),
    .Y(_109_));
 sky130_fd_sc_hd__nand2_1 _377_ (.A(_231_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__o21ai_1 _378_ (.A1(_229_),
    .A2(_109_),
    .B1(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_1 _379_ (.A1(_033_),
    .A2(_111_),
    .B1(_195_),
    .Y(_112_));
 sky130_fd_sc_hd__xnor2_1 _380_ (.A(_194_),
    .B(_112_),
    .Y(net68));
 sky130_fd_sc_hd__nor2_1 _381_ (.A(net2),
    .B(net34),
    .Y(_113_));
 sky130_fd_sc_hd__nor2_1 _382_ (.A(_113_),
    .B(_112_),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _383_ (.A(_193_),
    .B(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__xnor2_1 _384_ (.A(_192_),
    .B(_115_),
    .Y(net69));
 sky130_fd_sc_hd__mux2i_2 _385_ (.A0(_036_),
    .A1(_058_),
    .S(_109_),
    .Y(_116_));
 sky130_fd_sc_hd__xor2_1 _386_ (.A(_236_),
    .B(_116_),
    .X(net70));
 sky130_fd_sc_hd__inv_1 _387_ (.A(_235_),
    .Y(_117_));
 sky130_fd_sc_hd__mux2i_1 _388_ (.A0(_237_),
    .A1(_117_),
    .S(_116_),
    .Y(_118_));
 sky130_fd_sc_hd__xnor2_1 _389_ (.A(_202_),
    .B(_118_),
    .Y(net71));
 sky130_fd_sc_hd__nor2_1 _390_ (.A(net5),
    .B(net37),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_119_),
    .B(_118_),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_1 _392_ (.A(_201_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__xnor2_1 _393_ (.A(_200_),
    .B(_121_),
    .Y(net72));
 sky130_fd_sc_hd__o21bai_1 _394_ (.A1(_039_),
    .A2(_121_),
    .B1_N(_199_),
    .Y(_122_));
 sky130_fd_sc_hd__xor2_1 _395_ (.A(_198_),
    .B(_122_),
    .X(net73));
 sky130_fd_sc_hd__xor2_1 _396_ (.A(_248_),
    .B(_064_),
    .X(net74));
 sky130_fd_sc_hd__nand3_1 _397_ (.A(_247_),
    .B(_052_),
    .C(_062_),
    .Y(_123_));
 sky130_fd_sc_hd__o21ai_1 _398_ (.A1(_153_),
    .A2(_064_),
    .B1(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__xnor2_1 _399_ (.A(_208_),
    .B(_124_),
    .Y(net75));
 sky130_fd_sc_hd__o21a_1 _400_ (.A1(_002_),
    .A2(_124_),
    .B1(_001_),
    .X(_125_));
 sky130_fd_sc_hd__xnor2_1 _401_ (.A(_206_),
    .B(_125_),
    .Y(net76));
 sky130_fd_sc_hd__nor2_1 _402_ (.A(_004_),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _403_ (.A(_205_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(_204_),
    .B(_127_),
    .Y(net77));
 sky130_fd_sc_hd__and2_0 _405_ (.A(_016_),
    .B(_017_),
    .X(_128_));
 sky130_fd_sc_hd__xnor2_1 _406_ (.A(_184_),
    .B(_128_),
    .Y(net78));
 sky130_fd_sc_hd__xor2_1 _407_ (.A(_158_),
    .B(_087_),
    .X(net79));
 sky130_fd_sc_hd__inv_1 _408_ (.A(_157_),
    .Y(_129_));
 sky130_fd_sc_hd__mux2i_1 _409_ (.A0(_159_),
    .A1(_129_),
    .S(_087_),
    .Y(_130_));
 sky130_fd_sc_hd__xnor2_1 _410_ (.A(_214_),
    .B(_130_),
    .Y(net80));
 sky130_fd_sc_hd__o21bai_1 _411_ (.A1(_008_),
    .A2(_130_),
    .B1_N(_213_),
    .Y(_131_));
 sky130_fd_sc_hd__xor2_1 _412_ (.A(_212_),
    .B(_131_),
    .X(net81));
 sky130_fd_sc_hd__xnor2_1 _413_ (.A(_210_),
    .B(_074_),
    .Y(net82));
 sky130_fd_sc_hd__a31oi_4 _414_ (.A1(_065_),
    .A2(_073_),
    .A3(_083_),
    .B1(_209_),
    .Y(_132_));
 sky130_fd_sc_hd__xnor2_1 _415_ (.A(_164_),
    .B(_132_),
    .Y(net83));
 sky130_fd_sc_hd__inv_1 _416_ (.A(_163_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2i_2 _417_ (.A0(_133_),
    .A1(_165_),
    .S(_132_),
    .Y(_134_));
 sky130_fd_sc_hd__xnor2_1 _418_ (.A(_220_),
    .B(_134_),
    .Y(net84));
 sky130_fd_sc_hd__o21ba_1 _419_ (.A1(_075_),
    .A2(_134_),
    .B1_N(_219_),
    .X(_135_));
 sky130_fd_sc_hd__xnor2_1 _420_ (.A(_218_),
    .B(_135_),
    .Y(net85));
 sky130_fd_sc_hd__mux2i_1 _421_ (.A0(_078_),
    .A1(_091_),
    .S(_132_),
    .Y(_136_));
 sky130_fd_sc_hd__xor2_1 _422_ (.A(_216_),
    .B(_136_),
    .X(net86));
 sky130_fd_sc_hd__mux2i_1 _423_ (.A0(_080_),
    .A1(_097_),
    .S(_132_),
    .Y(_137_));
 sky130_fd_sc_hd__xor2_1 _424_ (.A(_170_),
    .B(_137_),
    .X(net87));
 sky130_fd_sc_hd__xor2_1 _425_ (.A(_226_),
    .B(_104_),
    .X(net88));
 sky130_fd_sc_hd__nor2_1 _426_ (.A(net12),
    .B(net44),
    .Y(_138_));
 sky130_fd_sc_hd__nor2_1 _427_ (.A(_128_),
    .B(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__nor2_1 _428_ (.A(_183_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_1 _429_ (.A(_182_),
    .B(_140_),
    .Y(net89));
 sky130_fd_sc_hd__xnor2_1 _430_ (.A(_224_),
    .B(_105_),
    .Y(net90));
 sky130_fd_sc_hd__o2111ai_1 _431_ (.A1(net24),
    .A2(net56),
    .B1(_222_),
    .C1(_000_),
    .D1(_104_),
    .Y(_141_));
 sky130_fd_sc_hd__or4_1 _432_ (.A(_222_),
    .B(_223_),
    .C(_225_),
    .D(_104_),
    .X(_142_));
 sky130_fd_sc_hd__o211ai_1 _433_ (.A1(net24),
    .A2(net56),
    .B1(_222_),
    .C1(_225_),
    .Y(_143_));
 sky130_fd_sc_hd__o41ai_1 _434_ (.A1(net24),
    .A2(net56),
    .A3(_222_),
    .A4(_223_),
    .B1(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__nor4_1 _435_ (.A(_222_),
    .B(_223_),
    .C(_225_),
    .D(_000_),
    .Y(_145_));
 sky130_fd_sc_hd__a211oi_1 _436_ (.A1(_222_),
    .A2(_223_),
    .B1(_144_),
    .C1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__and3_1 _437_ (.A(_141_),
    .B(_142_),
    .C(_146_),
    .X(net91));
 sky130_fd_sc_hd__xor2_1 _438_ (.A(_180_),
    .B(_021_),
    .X(net92));
 sky130_fd_sc_hd__xnor2_1 _439_ (.A(_176_),
    .B(_022_),
    .Y(net93));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(_177_),
    .B(_022_),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_1 _441_ (.A1(_175_),
    .A2(_022_),
    .B1(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__xor2_1 _442_ (.A(_190_),
    .B(_148_),
    .X(net94));
 sky130_fd_sc_hd__or2_0 _443_ (.A(net28),
    .B(net60),
    .X(_149_));
 sky130_fd_sc_hd__a21oi_1 _444_ (.A1(_149_),
    .A2(_148_),
    .B1(_189_),
    .Y(_150_));
 sky130_fd_sc_hd__xnor2_1 _445_ (.A(_188_),
    .B(_150_),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _446_ (.A(_025_),
    .Y(_151_));
 sky130_fd_sc_hd__a21oi_1 _447_ (.A1(_151_),
    .A2(_148_),
    .B1(_024_),
    .Y(_152_));
 sky130_fd_sc_hd__xnor2_1 _448_ (.A(_186_),
    .B(_152_),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_1 _449_ (.A(_230_),
    .B(_109_),
    .Y(net97));
 sky130_fd_sc_hd__xor2_1 _450_ (.A(_196_),
    .B(_111_),
    .X(net98));
 sky130_fd_sc_hd__ha_1 _451_ (.A(net8),
    .B(net40),
    .COUT(_153_),
    .SUM(_154_));
 sky130_fd_sc_hd__ha_1 _452_ (.A(_155_),
    .B(_156_),
    .COUT(_157_),
    .SUM(_158_));
 sky130_fd_sc_hd__ha_1 _453_ (.A(net13),
    .B(net45),
    .COUT(_159_),
    .SUM(_160_));
 sky130_fd_sc_hd__ha_1 _454_ (.A(_161_),
    .B(_162_),
    .COUT(_163_),
    .SUM(_164_));
 sky130_fd_sc_hd__ha_1 _455_ (.A(net17),
    .B(net49),
    .COUT(_165_),
    .SUM(_166_));
 sky130_fd_sc_hd__ha_1 _456_ (.A(_167_),
    .B(_168_),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__ha_1 _457_ (.A(net21),
    .B(net53),
    .COUT(_171_),
    .SUM(_172_));
 sky130_fd_sc_hd__ha_1 _458_ (.A(_173_),
    .B(_174_),
    .COUT(_175_),
    .SUM(_176_));
 sky130_fd_sc_hd__ha_1 _459_ (.A(net27),
    .B(net59),
    .COUT(_177_),
    .SUM(_178_));
 sky130_fd_sc_hd__ha_1 _460_ (.A(net26),
    .B(net58),
    .COUT(_179_),
    .SUM(_180_));
 sky130_fd_sc_hd__ha_1 _461_ (.A(net23),
    .B(net55),
    .COUT(_181_),
    .SUM(_182_));
 sky130_fd_sc_hd__ha_1 _462_ (.A(net12),
    .B(net44),
    .COUT(_183_),
    .SUM(_184_));
 sky130_fd_sc_hd__ha_1 _463_ (.A(net30),
    .B(net62),
    .COUT(_185_),
    .SUM(_186_));
 sky130_fd_sc_hd__ha_1 _464_ (.A(net29),
    .B(net61),
    .COUT(_187_),
    .SUM(_188_));
 sky130_fd_sc_hd__ha_1 _465_ (.A(net28),
    .B(net60),
    .COUT(_189_),
    .SUM(_190_));
 sky130_fd_sc_hd__ha_1 _466_ (.A(net3),
    .B(net35),
    .COUT(_191_),
    .SUM(_192_));
 sky130_fd_sc_hd__ha_1 _467_ (.A(net2),
    .B(net34),
    .COUT(_193_),
    .SUM(_194_));
 sky130_fd_sc_hd__ha_1 _468_ (.A(net32),
    .B(net64),
    .COUT(_195_),
    .SUM(_196_));
 sky130_fd_sc_hd__ha_1 _469_ (.A(net7),
    .B(net39),
    .COUT(_197_),
    .SUM(_198_));
 sky130_fd_sc_hd__ha_1 _470_ (.A(net6),
    .B(net38),
    .COUT(_199_),
    .SUM(_200_));
 sky130_fd_sc_hd__ha_1 _471_ (.A(net5),
    .B(net37),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__ha_1 _472_ (.A(net11),
    .B(net43),
    .COUT(_203_),
    .SUM(_204_));
 sky130_fd_sc_hd__ha_1 _473_ (.A(net10),
    .B(net42),
    .COUT(_205_),
    .SUM(_206_));
 sky130_fd_sc_hd__ha_1 _474_ (.A(net9),
    .B(net41),
    .COUT(_207_),
    .SUM(_208_));
 sky130_fd_sc_hd__ha_2 _475_ (.A(net16),
    .B(net48),
    .COUT(_209_),
    .SUM(_210_));
 sky130_fd_sc_hd__ha_1 _476_ (.A(net15),
    .B(net47),
    .COUT(_211_),
    .SUM(_212_));
 sky130_fd_sc_hd__ha_1 _477_ (.A(net14),
    .B(net46),
    .COUT(_213_),
    .SUM(_214_));
 sky130_fd_sc_hd__ha_1 _478_ (.A(net20),
    .B(net52),
    .COUT(_215_),
    .SUM(_216_));
 sky130_fd_sc_hd__ha_1 _479_ (.A(net19),
    .B(net51),
    .COUT(_217_),
    .SUM(_218_));
 sky130_fd_sc_hd__ha_1 _480_ (.A(net18),
    .B(net50),
    .COUT(_219_),
    .SUM(_220_));
 sky130_fd_sc_hd__ha_1 _481_ (.A(net25),
    .B(net57),
    .COUT(_221_),
    .SUM(_222_));
 sky130_fd_sc_hd__ha_1 _482_ (.A(net24),
    .B(net56),
    .COUT(_223_),
    .SUM(_224_));
 sky130_fd_sc_hd__ha_1 _483_ (.A(net22),
    .B(net54),
    .COUT(_225_),
    .SUM(_226_));
 sky130_fd_sc_hd__ha_1 _484_ (.A(_227_),
    .B(_228_),
    .COUT(_229_),
    .SUM(_230_));
 sky130_fd_sc_hd__ha_1 _485_ (.A(net31),
    .B(net63),
    .COUT(_231_),
    .SUM(_232_));
 sky130_fd_sc_hd__ha_1 _486_ (.A(_233_),
    .B(_234_),
    .COUT(_235_),
    .SUM(_236_));
 sky130_fd_sc_hd__ha_1 _487_ (.A(net4),
    .B(net36),
    .COUT(_237_),
    .SUM(_238_));
 sky130_fd_sc_hd__ha_1 _488_ (.A(_239_),
    .B(_240_),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__ha_1 _489_ (.A(net1),
    .B(net33),
    .COUT(_243_),
    .SUM(_244_));
 sky130_fd_sc_hd__ha_1 _490_ (.A(_245_),
    .B(_246_),
    .COUT(_247_),
    .SUM(_248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_43 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(sum[9]));
 sky130_fd_sc_hd__fill_2 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
endmodule
