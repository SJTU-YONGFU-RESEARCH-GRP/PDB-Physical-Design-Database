module barrel_shifter (rotate,
    shift_direction,
    data_in,
    data_out,
    shift_amount);
 input rotate;
 input shift_direction;
 input [31:0] data_in;
 output [31:0] data_out;
 input [4:0] shift_amount;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0812_ (.I(shift_amount[0]),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _0813_ (.I(_0641_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0814_ (.I(_0651_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0815_ (.I(_0662_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0816_ (.I(_0672_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0817_ (.I(net34),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _0818_ (.I(_0692_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0819_ (.I(net35),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _0820_ (.I(_0810_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _0821_ (.A1(net36),
    .A2(_0711_),
    .A3(_0721_),
    .B(net37),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0822_ (.A1(net37),
    .A2(net36),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _0823_ (.A1(_0711_),
    .A2(_0721_),
    .A3(_0742_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _0824_ (.I(_0641_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0825_ (.I(net34),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0826_ (.A1(_0711_),
    .A2(_0762_),
    .A3(_0772_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _0827_ (.A1(_0782_),
    .A2(_0742_),
    .B(net33),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0828_ (.A1(_0732_),
    .A2(_0752_),
    .B(_0792_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0829_ (.I(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0830_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0831_ (.I(net5),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0832_ (.I(_0811_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0833_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0834_ (.I0(_0803_),
    .I1(net7),
    .S(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0835_ (.I0(net4),
    .I1(net6),
    .S(_0804_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0836_ (.I(_0651_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0837_ (.I(_0000_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0838_ (.I0(_0806_),
    .I1(_0807_),
    .S(_0001_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0839_ (.I(net32),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0840_ (.I(net3),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0841_ (.I0(_0003_),
    .I1(_0004_),
    .S(_0805_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0842_ (.I(net31),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0843_ (.I(_0804_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0844_ (.I0(_0006_),
    .I1(net2),
    .S(_0007_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0845_ (.I0(_0005_),
    .I1(_0008_),
    .S(_0001_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _0846_ (.A1(net35),
    .A2(_0810_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0847_ (.I(_0010_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0848_ (.I(_0011_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0849_ (.I0(_0002_),
    .I1(_0009_),
    .S(_0012_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0850_ (.I(net28),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0851_ (.I(net30),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0852_ (.I(_0007_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0853_ (.I0(_0014_),
    .I1(_0015_),
    .S(_0016_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0854_ (.I(net27),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0855_ (.I(net29),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0856_ (.I0(_0018_),
    .I1(_0019_),
    .S(_0007_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0857_ (.I(net26),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0858_ (.I0(net12),
    .I1(_0021_),
    .S(_0016_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0859_ (.I(_0804_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0860_ (.I(_0023_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0861_ (.I0(net1),
    .I1(net23),
    .S(_0024_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0862_ (.I(_0010_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0863_ (.I(_0026_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0864_ (.I(_0027_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0865_ (.I0(_0017_),
    .I1(_0020_),
    .I2(_0022_),
    .I3(_0025_),
    .S0(_0808_),
    .S1(_0028_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0866_ (.I(net34),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0867_ (.A1(net36),
    .A2(_0711_),
    .A3(_0641_),
    .A4(_0030_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _0868_ (.A1(_0711_),
    .A2(_0641_),
    .A3(_0030_),
    .B(net36),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0869_ (.A1(_0031_),
    .A2(_0032_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0870_ (.I(_0033_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0871_ (.I(_0034_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0872_ (.I0(_0013_),
    .I1(_0029_),
    .S(_0035_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0873_ (.I(_0651_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _0874_ (.A1(net37),
    .A2(net36),
    .A3(net35),
    .A4(net34),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0875_ (.I(net33),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0876_ (.A1(_0037_),
    .A2(_0038_),
    .B(_0039_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0877_ (.A1(_0040_),
    .A2(_0732_),
    .A3(_0752_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0878_ (.I(_0041_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0879_ (.I(net21),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0880_ (.I0(_0043_),
    .I1(net22),
    .I2(net24),
    .I3(net25),
    .S0(_0641_),
    .S1(_0023_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0881_ (.I(net18),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0882_ (.I(net19),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0883_ (.I(_0804_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0884_ (.I0(net17),
    .I1(_0045_),
    .I2(_0046_),
    .I3(net20),
    .S0(_0762_),
    .S1(_0047_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0885_ (.I0(_0044_),
    .I1(_0048_),
    .S(_0026_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0886_ (.I0(net13),
    .I1(net14),
    .I2(net15),
    .I3(net16),
    .S0(_0762_),
    .S1(_0047_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0887_ (.I(net9),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0888_ (.I0(net8),
    .I1(_0051_),
    .I2(net10),
    .I3(net11),
    .S0(_0641_),
    .S1(_0047_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0889_ (.I0(_0050_),
    .I1(_0052_),
    .S(_0026_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0890_ (.I0(_0049_),
    .I1(_0053_),
    .S(_0033_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0891_ (.A1(_0802_),
    .A2(_0036_),
    .B1(_0042_),
    .B2(_0054_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0892_ (.A1(net1),
    .A2(_0000_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _0893_ (.I(net38),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0894_ (.I(_0057_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0895_ (.I(_0058_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0896_ (.A1(_0056_),
    .A2(_0038_),
    .B(_0059_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _0897_ (.I(_0023_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0898_ (.I(net36),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _0899_ (.A1(_0062_),
    .A2(_0782_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0900_ (.A1(_0810_),
    .A2(_0063_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0901_ (.I(_0711_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0902_ (.A1(_0065_),
    .A2(_0721_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0903_ (.I(_0641_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _0904_ (.A1(_0067_),
    .A2(_0692_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0905_ (.A1(_0065_),
    .A2(_0721_),
    .A3(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _0906_ (.A1(_0066_),
    .A2(_0069_),
    .B(_0062_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0907_ (.A1(_0064_),
    .A2(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _0908_ (.A1(_0061_),
    .A2(_0071_),
    .A3(_0801_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0909_ (.I(net38),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0910_ (.I(_0073_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0911_ (.I0(net18),
    .I1(net20),
    .S(_0030_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0912_ (.I0(net17),
    .I1(_0046_),
    .S(_0772_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0913_ (.I0(_0075_),
    .I1(_0076_),
    .S(_0037_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0914_ (.I0(net22),
    .I1(net25),
    .S(_0030_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0915_ (.I0(net21),
    .I1(net24),
    .S(_0030_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _0916_ (.I0(_0078_),
    .I1(_0079_),
    .S(_0651_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _0917_ (.I0(_0077_),
    .I1(_0080_),
    .S(_0065_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0918_ (.I(net13),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0919_ (.I(net14),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0920_ (.I(net15),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0921_ (.I(net16),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0922_ (.I(_0641_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0923_ (.I(_0692_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0924_ (.I0(_0082_),
    .I1(_0083_),
    .I2(_0084_),
    .I3(_0085_),
    .S0(_0086_),
    .S1(_0087_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0925_ (.I(net8),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0926_ (.I(net10),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0927_ (.I(net11),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0928_ (.I0(_0089_),
    .I1(_0051_),
    .I2(_0090_),
    .I3(_0091_),
    .S0(_0086_),
    .S1(_0087_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _0929_ (.I(_0711_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0930_ (.I(_0093_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0931_ (.I0(_0088_),
    .I1(_0092_),
    .S(_0094_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _0932_ (.I(_0062_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0933_ (.I0(_0081_),
    .I1(_0095_),
    .S(_0096_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0934_ (.I(net4),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0935_ (.I(net6),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0936_ (.I(_0641_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0937_ (.I0(_0098_),
    .I1(_0803_),
    .I2(_0099_),
    .I3(net7),
    .S0(_0100_),
    .S1(_0087_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0938_ (.I(net2),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0939_ (.I0(_0006_),
    .I1(_0003_),
    .I2(_0102_),
    .I3(_0004_),
    .S0(_0100_),
    .S1(_0087_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0940_ (.I0(_0101_),
    .I1(_0103_),
    .S(_0094_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0941_ (.I(_0692_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0942_ (.I0(_0018_),
    .I1(_0014_),
    .I2(_0019_),
    .I3(_0015_),
    .S0(_0100_),
    .S1(_0105_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0943_ (.I(_0762_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0944_ (.I0(net1),
    .I1(net12),
    .I2(net23),
    .I3(_0021_),
    .S0(_0107_),
    .S1(_0105_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0945_ (.I(_0093_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0946_ (.I0(_0106_),
    .I1(_0108_),
    .S(_0109_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0947_ (.I(_0096_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0948_ (.I0(_0104_),
    .I1(_0110_),
    .S(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0949_ (.I(net37),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0950_ (.I(_0113_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0951_ (.I0(_0097_),
    .I1(_0112_),
    .S(_0114_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _0952_ (.A1(_0056_),
    .A2(_0072_),
    .B(_0074_),
    .C(_0115_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0953_ (.A1(_0055_),
    .A2(_0060_),
    .B(_0116_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _0954_ (.I0(net24),
    .I1(net25),
    .S(_0641_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0955_ (.A1(_0061_),
    .A2(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0956_ (.I0(_0046_),
    .I1(net20),
    .I2(_0043_),
    .I3(net22),
    .S0(_0100_),
    .S1(_0024_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0957_ (.I0(_0118_),
    .I1(_0119_),
    .S(_0027_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0958_ (.I(_0033_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0959_ (.A1(_0732_),
    .A2(_0752_),
    .A3(_0121_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0960_ (.A1(_0732_),
    .A2(_0752_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _0961_ (.I0(_0090_),
    .I1(_0091_),
    .I2(_0082_),
    .I3(_0083_),
    .S0(_0100_),
    .S1(_0024_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0962_ (.I0(net3),
    .I1(net5),
    .S(_0804_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0963_ (.I0(_0102_),
    .I1(_0098_),
    .S(_0805_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0964_ (.I(_0651_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0965_ (.I0(_0125_),
    .I1(_0126_),
    .S(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0966_ (.I0(_0124_),
    .I1(_0128_),
    .S(_0033_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0967_ (.A1(_0123_),
    .A2(_0028_),
    .A3(_0129_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0968_ (.A1(_0120_),
    .A2(_0122_),
    .B(_0130_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _0969_ (.I(_0114_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0970_ (.I(_0065_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0971_ (.I(_0021_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0972_ (.I(_0018_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0973_ (.I(_0014_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0974_ (.I(_0019_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0975_ (.I0(_0134_),
    .I1(_0135_),
    .I2(_0136_),
    .I3(_0137_),
    .S0(_0127_),
    .S1(_0809_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0976_ (.I(net34),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0977_ (.I(_0139_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0978_ (.I0(_0102_),
    .I1(_0003_),
    .I2(_0006_),
    .I3(_0015_),
    .S0(_0086_),
    .S1(_0140_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0979_ (.A1(_0133_),
    .A2(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0980_ (.A1(_0133_),
    .A2(_0138_),
    .B(_0142_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0981_ (.I0(net23),
    .I1(net1),
    .S(_0030_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0982_ (.A1(net12),
    .A2(_0107_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _0983_ (.A1(_0672_),
    .A2(_0144_),
    .B1(_0145_),
    .B2(_0809_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0984_ (.A1(_0133_),
    .A2(_0146_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0985_ (.I0(_0143_),
    .I1(_0147_),
    .S(_0062_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0986_ (.A1(_0132_),
    .A2(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _0987_ (.A1(_0711_),
    .A2(_0810_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0988_ (.I(_0150_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0989_ (.I(_0151_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _0990_ (.I(net17),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _0991_ (.I0(_0084_),
    .I1(_0085_),
    .I2(_0153_),
    .I3(_0045_),
    .S0(_0067_),
    .S1(_0016_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0992_ (.I0(net7),
    .I1(net9),
    .S(_0804_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0993_ (.I0(_0099_),
    .I1(_0089_),
    .S(_0007_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0994_ (.I0(_0155_),
    .I1(_0156_),
    .S(_0662_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0995_ (.I0(_0154_),
    .I1(_0157_),
    .S(_0121_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0996_ (.A1(_0800_),
    .A2(_0152_),
    .A3(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0997_ (.A1(_0058_),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _0998_ (.A1(_0792_),
    .A2(_0131_),
    .B(_0149_),
    .C(_0160_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0999_ (.A1(_0040_),
    .A2(_0123_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1000_ (.I0(net23),
    .I1(net1),
    .S(_0023_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1001_ (.A1(_0001_),
    .A2(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1002_ (.A1(_0061_),
    .A2(_0145_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1003_ (.A1(_0164_),
    .A2(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1004_ (.A1(_0031_),
    .A2(_0032_),
    .A3(_0026_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1005_ (.I0(net2),
    .I1(_0006_),
    .S(_0007_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1006_ (.I0(_0019_),
    .I1(_0018_),
    .S(_0047_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1007_ (.I0(_0168_),
    .I1(_0169_),
    .S(_0150_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1008_ (.I0(_0014_),
    .I1(_0021_),
    .S(_0023_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1009_ (.I0(_0003_),
    .I1(_0015_),
    .S(_0805_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1010_ (.I0(_0171_),
    .I1(_0172_),
    .S(_0026_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1011_ (.I(_0762_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1012_ (.I(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1013_ (.I0(_0170_),
    .I1(_0173_),
    .S(_0175_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1014_ (.I(_0121_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1015_ (.A1(_0166_),
    .A2(_0167_),
    .B1(_0176_),
    .B2(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1016_ (.I0(_0084_),
    .I1(_0085_),
    .I2(_0153_),
    .I3(_0045_),
    .S0(_0762_),
    .S1(_0692_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1017_ (.I0(_0090_),
    .I1(_0091_),
    .I2(_0082_),
    .I3(_0083_),
    .S0(_0762_),
    .S1(_0692_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1018_ (.I0(_0179_),
    .I1(_0180_),
    .S(_0093_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1019_ (.I0(_0099_),
    .I1(net7),
    .I2(_0089_),
    .I3(_0051_),
    .S0(_0762_),
    .S1(_0140_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1020_ (.I0(_0102_),
    .I1(_0004_),
    .I2(_0098_),
    .I3(_0803_),
    .S0(_0762_),
    .S1(_0140_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1021_ (.I0(_0182_),
    .I1(_0183_),
    .S(_0093_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1022_ (.I(_0096_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1023_ (.I0(_0181_),
    .I1(_0184_),
    .S(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1024_ (.I0(net19),
    .I1(net21),
    .S(_0030_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1025_ (.I0(net20),
    .I1(net22),
    .S(_0030_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1026_ (.I0(_0187_),
    .I1(_0188_),
    .S(_0067_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1027_ (.A1(_0809_),
    .A2(_0117_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1028_ (.I0(_0189_),
    .I1(_0190_),
    .S(_0065_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1029_ (.A1(net37),
    .A2(_0096_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1030_ (.I(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1031_ (.A1(_0132_),
    .A2(_0186_),
    .B1(_0191_),
    .B2(_0193_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1032_ (.I(_0058_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1033_ (.A1(_0162_),
    .A2(_0178_),
    .B(_0194_),
    .C(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1034_ (.A1(_0161_),
    .A2(_0196_),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1035_ (.I(_0132_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1036_ (.I0(net29),
    .I1(_0018_),
    .S(_0772_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1037_ (.I0(net30),
    .I1(net28),
    .S(_0030_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1038_ (.I0(_0198_),
    .I1(_0199_),
    .S(_0037_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1039_ (.I0(_0004_),
    .I1(_0102_),
    .I2(_0003_),
    .I3(_0006_),
    .S0(_0086_),
    .S1(_0087_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1040_ (.I0(_0200_),
    .I1(_0201_),
    .S(_0094_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1041_ (.I(_0093_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1042_ (.I0(net26),
    .I1(net12),
    .S(_0030_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _1043_ (.I0(_0144_),
    .I1(_0204_),
    .S(_0651_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1044_ (.A1(_0203_),
    .A2(_0205_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1045_ (.I0(_0202_),
    .I1(_0206_),
    .S(_0062_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1046_ (.A1(_0031_),
    .A2(_0032_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1047_ (.I(_0208_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1048_ (.A1(_0801_),
    .A2(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1049_ (.I0(_0085_),
    .I1(_0153_),
    .I2(_0045_),
    .I3(_0046_),
    .S0(_0067_),
    .S1(_0016_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1050_ (.I0(_0091_),
    .I1(_0082_),
    .I2(_0083_),
    .I3(_0084_),
    .S0(_0067_),
    .S1(_0016_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1051_ (.I0(_0211_),
    .I1(_0212_),
    .S(_0026_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1052_ (.A1(_0197_),
    .A2(_0207_),
    .B1(_0210_),
    .B2(_0213_),
    .C(_0195_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1053_ (.I(_0040_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1054_ (.A1(_0127_),
    .A2(net25),
    .A3(_0061_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1055_ (.I0(net20),
    .I1(_0043_),
    .I2(net22),
    .I3(net24),
    .S0(_0067_),
    .S1(_0016_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1056_ (.I0(_0216_),
    .I1(_0217_),
    .S(_0026_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1057_ (.I0(_0089_),
    .I1(net10),
    .S(_0007_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1058_ (.I0(_0219_),
    .I1(_0155_),
    .S(_0037_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1059_ (.I0(_0807_),
    .I1(_0125_),
    .S(_0037_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1060_ (.I0(_0220_),
    .I1(_0221_),
    .S(_0011_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1061_ (.I(_0123_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1062_ (.I0(_0218_),
    .I1(_0222_),
    .S(_0223_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1063_ (.A1(_0215_),
    .A2(_0035_),
    .A3(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1064_ (.I0(_0085_),
    .I1(_0153_),
    .I2(_0045_),
    .I3(_0046_),
    .S0(_0174_),
    .S1(_0105_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1065_ (.I0(_0091_),
    .I1(_0082_),
    .I2(_0083_),
    .I3(_0084_),
    .S0(_0100_),
    .S1(_0105_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1066_ (.I(_0093_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1067_ (.I(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1068_ (.I0(_0226_),
    .I1(_0227_),
    .S(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1069_ (.I0(net7),
    .I1(_0089_),
    .I2(_0051_),
    .I3(_0090_),
    .S0(_0100_),
    .S1(_0087_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1070_ (.I0(_0004_),
    .I1(_0098_),
    .I2(_0803_),
    .I3(_0099_),
    .S0(_0107_),
    .S1(_0105_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1071_ (.I0(_0231_),
    .I1(_0232_),
    .S(_0203_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1072_ (.I(_0096_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1073_ (.I(_0234_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1074_ (.I0(_0230_),
    .I1(_0233_),
    .S(_0235_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1075_ (.A1(_0809_),
    .A2(net25),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1076_ (.I0(_0188_),
    .I1(_0237_),
    .S(_0133_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1077_ (.A1(_0203_),
    .A2(_0079_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _1078_ (.I0(_0238_),
    .I1(_0239_),
    .S(_0175_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1079_ (.A1(_0197_),
    .A2(_0236_),
    .B1(_0240_),
    .B2(_0193_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1080_ (.I0(_0015_),
    .I1(_0014_),
    .S(_0047_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1081_ (.I0(_0169_),
    .I1(_0242_),
    .S(_0000_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1082_ (.I0(net3),
    .I1(_0003_),
    .S(_0007_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1083_ (.I0(_0168_),
    .I1(_0244_),
    .S(_0127_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1084_ (.I0(_0243_),
    .I1(_0245_),
    .S(_0027_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1085_ (.I0(_0021_),
    .I1(net12),
    .S(_0805_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1086_ (.I0(_0163_),
    .I1(_0247_),
    .S(_0000_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1087_ (.A1(_0012_),
    .A2(_0248_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1088_ (.I0(_0246_),
    .I1(_0249_),
    .S(_0209_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1089_ (.A1(_0802_),
    .A2(_0250_),
    .B(_0074_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1090_ (.A1(_0214_),
    .A2(_0225_),
    .B1(_0241_),
    .B2(_0251_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _1091_ (.I(_0801_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1092_ (.A1(net1),
    .A2(_0000_),
    .A3(_0061_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1093_ (.A1(_0711_),
    .A2(_0692_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1094_ (.A1(_0062_),
    .A2(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1095_ (.A1(_0151_),
    .A2(_0253_),
    .A3(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1096_ (.I0(_0018_),
    .I1(net23),
    .S(_0805_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1097_ (.I0(_0247_),
    .I1(_0257_),
    .S(_0000_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1098_ (.A1(_0027_),
    .A2(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1099_ (.I0(_0006_),
    .I1(_0019_),
    .S(_0023_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1100_ (.I0(_0098_),
    .I1(_0102_),
    .S(_0047_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1101_ (.I0(_0242_),
    .I1(_0244_),
    .I2(_0260_),
    .I3(_0261_),
    .S0(_0011_),
    .S1(_0001_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1102_ (.I0(_0259_),
    .I1(_0262_),
    .S(_0034_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1103_ (.A1(_0256_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1104_ (.A1(_0229_),
    .A2(_0193_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1105_ (.I(net38),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1106_ (.A1(_0252_),
    .A2(_0264_),
    .B1(_0265_),
    .B2(_0080_),
    .C(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1107_ (.I0(_0077_),
    .I1(_0088_),
    .S(_0229_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1108_ (.I0(_0092_),
    .I1(_0101_),
    .S(_0203_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1109_ (.I0(_0268_),
    .I1(_0269_),
    .S(_0235_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1110_ (.A1(_0197_),
    .A2(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1111_ (.A1(_0223_),
    .A2(_0209_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1112_ (.I0(_0048_),
    .I1(_0050_),
    .S(_0028_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1113_ (.A1(_0033_),
    .A2(_0044_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1114_ (.A1(_0732_),
    .A2(_0752_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1115_ (.I0(_0002_),
    .I1(_0274_),
    .S(_0275_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1116_ (.A1(_0028_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1117_ (.A1(_0152_),
    .A2(_0052_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1118_ (.I(_0275_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1119_ (.A1(_0035_),
    .A2(_0278_),
    .B(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _1120_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0277_),
    .B2(_0280_),
    .C(_0215_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1121_ (.A1(net1),
    .A2(_0068_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1122_ (.I0(net27),
    .I1(net23),
    .S(_0772_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1123_ (.I0(_0204_),
    .I1(_0283_),
    .S(_0037_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1124_ (.I0(_0282_),
    .I1(_0284_),
    .S(_0094_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1125_ (.I0(net31),
    .I1(_0019_),
    .S(_0772_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1126_ (.I0(_0199_),
    .I1(_0286_),
    .S(_0037_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1127_ (.I0(_0098_),
    .I1(_0004_),
    .I2(_0102_),
    .I3(_0003_),
    .S0(_0100_),
    .S1(_0087_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1128_ (.I0(_0287_),
    .I1(_0288_),
    .S(_0228_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1129_ (.I0(_0285_),
    .I1(_0289_),
    .S(_0234_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1130_ (.A1(_0197_),
    .A2(_0290_),
    .B(_0059_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1131_ (.A1(_0267_),
    .A2(_0271_),
    .B1(_0281_),
    .B2(_0291_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _1132_ (.I0(_0083_),
    .I1(_0084_),
    .I2(_0085_),
    .I3(_0153_),
    .S0(_0086_),
    .S1(_0024_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1133_ (.I0(_0045_),
    .I1(_0046_),
    .I2(net20),
    .I3(_0043_),
    .S0(_0086_),
    .S1(_0024_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1134_ (.I0(_0292_),
    .I1(_0293_),
    .S(_0151_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1135_ (.I0(_0806_),
    .I1(_0156_),
    .S(_0107_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1136_ (.I0(net22),
    .I1(net25),
    .S(_0047_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1137_ (.A1(_0174_),
    .A2(net24),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1138_ (.A1(_0672_),
    .A2(_0296_),
    .B1(_0297_),
    .B2(_0061_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1139_ (.I(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1140_ (.A1(_0223_),
    .A2(_0295_),
    .B1(_0299_),
    .B2(_0122_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _1141_ (.I0(_0051_),
    .I1(_0090_),
    .I2(_0091_),
    .I3(_0082_),
    .S0(_0067_),
    .S1(_0016_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1142_ (.A1(_0152_),
    .A2(_0301_),
    .B(_0209_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1143_ (.A1(_0152_),
    .A2(_0300_),
    .B1(_0302_),
    .B2(_0279_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1144_ (.A1(_0272_),
    .A2(_0294_),
    .B(_0303_),
    .C(_0215_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1145_ (.I0(_0014_),
    .I1(_0021_),
    .S(_0772_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1146_ (.I0(_0305_),
    .I1(_0283_),
    .S(_0107_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _1147_ (.I0(net12),
    .I1(net1),
    .S(_0762_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1148_ (.A1(_0809_),
    .A2(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1149_ (.I0(_0306_),
    .I1(_0308_),
    .S(_0065_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1150_ (.I0(net32),
    .I1(_0015_),
    .S(_0772_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1151_ (.I0(_0310_),
    .I1(_0286_),
    .S(_0107_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1152_ (.I0(_0803_),
    .I1(_0098_),
    .I2(_0004_),
    .I3(_0102_),
    .S0(_0067_),
    .S1(_0140_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1153_ (.I0(_0311_),
    .I1(_0312_),
    .S(_0094_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1154_ (.I0(_0309_),
    .I1(_0313_),
    .S(_0111_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1155_ (.A1(_0197_),
    .A2(_0314_),
    .B(_0059_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1156_ (.A1(_0061_),
    .A2(_0307_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1157_ (.I0(_0171_),
    .I1(_0257_),
    .S(_0174_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1158_ (.I0(_0316_),
    .I1(_0317_),
    .S(_0027_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1159_ (.I0(_0803_),
    .I1(_0004_),
    .S(_0023_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _1160_ (.I0(_0172_),
    .I1(_0260_),
    .I2(_0319_),
    .I3(_0261_),
    .S0(_0175_),
    .S1(_0012_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1161_ (.I0(_0318_),
    .I1(_0320_),
    .S(_0177_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _1162_ (.I0(_0051_),
    .I1(_0090_),
    .I2(_0091_),
    .I3(_0082_),
    .S0(_0086_),
    .S1(_0140_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1163_ (.I0(_0803_),
    .I1(_0099_),
    .I2(net7),
    .I3(_0089_),
    .S0(_0086_),
    .S1(_0087_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1164_ (.I0(_0322_),
    .I1(_0323_),
    .S(_0203_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1165_ (.A1(_0809_),
    .A2(net24),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1166_ (.I0(_0078_),
    .I1(_0325_),
    .S(_0175_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1167_ (.A1(_0229_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1168_ (.I(net37),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1169_ (.I0(_0324_),
    .I1(_0327_),
    .S(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1170_ (.I(_0062_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1171_ (.I0(_0083_),
    .I1(_0084_),
    .I2(_0085_),
    .I3(_0153_),
    .S0(_0086_),
    .S1(_0140_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1172_ (.I0(_0075_),
    .I1(_0187_),
    .S(_0174_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1173_ (.I0(_0331_),
    .I1(_0332_),
    .S(_0133_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1174_ (.A1(_0114_),
    .A2(_0330_),
    .A3(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1175_ (.A1(_0073_),
    .A2(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1176_ (.A1(_0252_),
    .A2(_0321_),
    .B1(_0329_),
    .B2(_0235_),
    .C(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1177_ (.A1(_0304_),
    .A2(_0315_),
    .B(_0336_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1178_ (.I(_0328_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1179_ (.I0(_0124_),
    .I1(_0157_),
    .S(_0011_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1180_ (.A1(_0275_),
    .A2(_0209_),
    .A3(_0338_),
    .B(_0040_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1181_ (.A1(_0065_),
    .A2(_0721_),
    .A3(_0068_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1182_ (.A1(_0328_),
    .A2(_0068_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1183_ (.A1(_0096_),
    .A2(_0093_),
    .A3(_0810_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1184_ (.A1(_0096_),
    .A2(_0340_),
    .B(_0341_),
    .C(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1185_ (.A1(_0118_),
    .A2(_0343_),
    .B(_0123_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1186_ (.I0(_0119_),
    .I1(_0154_),
    .S(_0011_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1187_ (.A1(_0275_),
    .A2(_0034_),
    .A3(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1188_ (.A1(_0339_),
    .A2(_0344_),
    .A3(_0346_),
    .B(_0073_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1189_ (.I0(_0169_),
    .I1(_0171_),
    .S(_0175_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1190_ (.A1(_0012_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1191_ (.A1(_0152_),
    .A2(_0166_),
    .B(_0349_),
    .C(_0177_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1192_ (.I0(_0099_),
    .I1(_0098_),
    .S(_0007_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1193_ (.I0(_0319_),
    .I1(_0351_),
    .S(_0000_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1194_ (.A1(_0064_),
    .A2(_0070_),
    .B(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1195_ (.I0(_0168_),
    .I1(_0172_),
    .S(_0174_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1196_ (.A1(_0711_),
    .A2(_0810_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1197_ (.A1(_0065_),
    .A2(_0810_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1198_ (.A1(_0068_),
    .A2(_0355_),
    .B(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1199_ (.A1(_0721_),
    .A2(_0063_),
    .B1(_0357_),
    .B2(_0062_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1200_ (.A1(_0354_),
    .A2(_0358_),
    .B(_0801_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1201_ (.A1(_0254_),
    .A2(_0192_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1202_ (.A1(_0117_),
    .A2(_0360_),
    .B(net38),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1203_ (.A1(_0350_),
    .A2(_0353_),
    .A3(_0359_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1204_ (.A1(_0347_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1205_ (.I0(_0179_),
    .I1(_0189_),
    .S(_0133_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1206_ (.I0(_0180_),
    .I1(_0182_),
    .S(_0228_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1207_ (.I0(_0364_),
    .I1(_0365_),
    .S(_0235_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1208_ (.A1(_0362_),
    .A2(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1209_ (.A1(_0339_),
    .A2(_0344_),
    .A3(_0346_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1210_ (.I0(_0138_),
    .I1(_0146_),
    .S(_0133_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1211_ (.I0(_0099_),
    .I1(_0803_),
    .I2(_0098_),
    .I3(_0004_),
    .S0(_0100_),
    .S1(_0087_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1212_ (.I0(_0141_),
    .I1(_0370_),
    .S(_0228_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1213_ (.I(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1214_ (.I0(_0369_),
    .I1(_0372_),
    .S(_0185_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1215_ (.A1(_0266_),
    .A2(_0368_),
    .A3(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1216_ (.A1(_0337_),
    .A2(_0363_),
    .B(_0367_),
    .C(_0374_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1217_ (.I0(_0211_),
    .I1(_0217_),
    .S(_0150_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1218_ (.A1(_0279_),
    .A2(_0177_),
    .A3(_0375_),
    .B(_0040_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1219_ (.A1(_0216_),
    .A2(_0343_),
    .B(_0223_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1220_ (.I0(_0212_),
    .I1(_0220_),
    .S(_0011_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1221_ (.A1(_0279_),
    .A2(_0209_),
    .A3(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _1222_ (.A1(_0376_),
    .A2(_0377_),
    .A3(_0379_),
    .B(_0073_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1223_ (.I0(_0243_),
    .I1(_0248_),
    .S(_0151_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1224_ (.A1(_0177_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1225_ (.I0(net7),
    .I1(_0803_),
    .S(_0007_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1226_ (.I0(_0351_),
    .I1(_0383_),
    .S(_0127_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1227_ (.A1(_0064_),
    .A2(_0070_),
    .B(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1228_ (.A1(_0245_),
    .A2(_0358_),
    .B(_0800_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1229_ (.A1(_0808_),
    .A2(net25),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1230_ (.A1(_0387_),
    .A2(_0360_),
    .B(net38),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _1231_ (.A1(_0382_),
    .A2(_0385_),
    .A3(_0386_),
    .B(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1232_ (.A1(_0380_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1233_ (.I0(_0200_),
    .I1(_0205_),
    .S(_0065_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1234_ (.I0(_0099_),
    .I1(net4),
    .S(_0772_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1235_ (.I0(net7),
    .I1(_0803_),
    .S(_0772_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1236_ (.I0(_0392_),
    .I1(_0393_),
    .S(_0037_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1237_ (.I0(_0201_),
    .I1(_0394_),
    .S(_0094_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1238_ (.I0(_0391_),
    .I1(_0395_),
    .S(_0111_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1239_ (.I0(_0079_),
    .I1(_0188_),
    .S(_0672_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1240_ (.I0(_0226_),
    .I1(_0397_),
    .S(_0133_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1241_ (.I0(_0227_),
    .I1(_0231_),
    .S(_0109_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1242_ (.I0(_0398_),
    .I1(_0399_),
    .S(_0185_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1243_ (.A1(_0380_),
    .A2(_0396_),
    .B1(_0389_),
    .B2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1244_ (.A1(_0337_),
    .A2(_0390_),
    .B(_0401_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1245_ (.I(_0073_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1246_ (.I0(_0257_),
    .I1(_0260_),
    .S(_0026_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1247_ (.A1(_0808_),
    .A2(_0031_),
    .A3(_0032_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1248_ (.I0(_0242_),
    .I1(_0247_),
    .S(_0150_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1249_ (.A1(_0330_),
    .A2(_0808_),
    .A3(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1250_ (.A1(_0403_),
    .A2(_0404_),
    .B(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1251_ (.I0(_0089_),
    .I1(_0099_),
    .S(_0023_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1252_ (.I0(_0383_),
    .I1(_0408_),
    .S(_0000_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1253_ (.A1(_0064_),
    .A2(_0070_),
    .B(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1254_ (.I0(_0244_),
    .I1(_0261_),
    .S(_0672_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1255_ (.A1(_0358_),
    .A2(_0411_),
    .B(_0800_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _1256_ (.A1(_0407_),
    .A2(_0410_),
    .A3(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1257_ (.A1(_0071_),
    .A2(_0042_),
    .A3(_0253_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1258_ (.A1(_0800_),
    .A2(_0054_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1259_ (.A1(_0056_),
    .A2(_0360_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1260_ (.A1(_0058_),
    .A2(_0415_),
    .A3(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1261_ (.A1(_0402_),
    .A2(_0413_),
    .A3(_0414_),
    .B(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1262_ (.I0(_0284_),
    .I1(_0287_),
    .S(_0094_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1263_ (.I0(_0089_),
    .I1(_0099_),
    .S(_0139_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1264_ (.I0(_0393_),
    .I1(_0420_),
    .S(_0662_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1265_ (.I0(_0288_),
    .I1(_0421_),
    .S(_0109_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1266_ (.I0(_0419_),
    .I1(_0422_),
    .S(_0235_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1267_ (.A1(_0417_),
    .A2(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _1268_ (.A1(_0074_),
    .A2(_0097_),
    .A3(_0413_),
    .A4(_0414_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1269_ (.A1(_0337_),
    .A2(_0418_),
    .B(_0424_),
    .C(_0425_),
    .ZN(net46));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1270_ (.A1(_0316_),
    .A2(_0343_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1271_ (.I0(_0173_),
    .I1(_0403_),
    .S(_0175_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1272_ (.A1(_0279_),
    .A2(_0177_),
    .A3(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1273_ (.A1(_0279_),
    .A2(_0426_),
    .B(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1274_ (.I0(_0261_),
    .I1(_0408_),
    .S(_0026_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1275_ (.I0(_0051_),
    .I1(net7),
    .S(_0047_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1276_ (.I0(_0319_),
    .I1(_0431_),
    .S(_0026_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1277_ (.I0(_0430_),
    .I1(_0432_),
    .S(_0001_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1278_ (.A1(_0279_),
    .A2(_0209_),
    .A3(_0433_),
    .B(_0040_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1279_ (.A1(_0058_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1280_ (.A1(_0150_),
    .A2(_0293_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1281_ (.A1(_0151_),
    .A2(_0298_),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1282_ (.A1(_0292_),
    .A2(_0358_),
    .B1(_0437_),
    .B2(_0177_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1283_ (.A1(_0064_),
    .A2(_0070_),
    .B(_0301_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1284_ (.A1(_0307_),
    .A2(_0360_),
    .B(_0057_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1285_ (.A1(_0162_),
    .A2(_0438_),
    .A3(_0439_),
    .B(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1286_ (.A1(_0402_),
    .A2(_0429_),
    .B(_0435_),
    .C(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1287_ (.I0(_0306_),
    .I1(_0311_),
    .S(_0203_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1288_ (.I0(_0051_),
    .I1(net7),
    .S(_0772_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1289_ (.I0(_0420_),
    .I1(_0444_),
    .S(_0037_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1290_ (.I0(_0312_),
    .I1(_0445_),
    .S(_0229_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1291_ (.I0(_0443_),
    .I1(_0446_),
    .S(_0235_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1292_ (.A1(_0441_),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1293_ (.A1(_0275_),
    .A2(_0209_),
    .A3(_0433_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1294_ (.A1(_0215_),
    .A2(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _1295_ (.I0(_0075_),
    .I1(_0078_),
    .I2(_0187_),
    .I3(_0325_),
    .S0(_0065_),
    .S1(_0174_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1296_ (.I0(_0331_),
    .I1(_0322_),
    .S(_0093_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1297_ (.I0(_0451_),
    .I1(_0452_),
    .S(_0111_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1298_ (.A1(_0429_),
    .A2(_0450_),
    .B(_0453_),
    .C(_0266_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1299_ (.A1(_0337_),
    .A2(_0442_),
    .B(_0448_),
    .C(_0454_),
    .ZN(net47));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1300_ (.I0(_0181_),
    .I1(_0191_),
    .S(_0062_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1301_ (.A1(_0071_),
    .A2(_0042_),
    .A3(_0166_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1302_ (.A1(_0197_),
    .A2(_0455_),
    .B(_0456_),
    .C(_0074_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1303_ (.I0(_0090_),
    .I1(_0089_),
    .S(_0805_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1304_ (.I0(_0351_),
    .I1(_0458_),
    .S(_0027_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1305_ (.I0(_0432_),
    .I1(_0459_),
    .S(_0808_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1306_ (.I0(_0176_),
    .I1(_0460_),
    .S(_0035_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1307_ (.A1(_0802_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1308_ (.I0(_0124_),
    .I1(_0154_),
    .S(_0151_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1309_ (.I0(_0120_),
    .I1(_0463_),
    .S(_0034_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1310_ (.I0(_0090_),
    .I1(_0089_),
    .S(_0139_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1311_ (.I0(_0444_),
    .I1(_0465_),
    .S(_0662_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1312_ (.I0(_0370_),
    .I1(_0466_),
    .S(_0109_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1313_ (.I0(_0143_),
    .I1(_0467_),
    .S(_0185_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1314_ (.A1(_0229_),
    .A2(_0193_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1315_ (.A1(_0146_),
    .A2(_0469_),
    .B(_0073_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1316_ (.A1(_0252_),
    .A2(_0464_),
    .B1(_0468_),
    .B2(_0132_),
    .C(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1317_ (.A1(_0457_),
    .A2(_0462_),
    .B(_0471_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1318_ (.I0(_0213_),
    .I1(_0218_),
    .S(_0208_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1319_ (.A1(_0205_),
    .A2(_0265_),
    .B1(_0472_),
    .B2(_0252_),
    .C(_0195_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1320_ (.I0(net11),
    .I1(_0051_),
    .S(_0139_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1321_ (.I0(_0465_),
    .I1(_0474_),
    .S(_0662_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1322_ (.I0(_0394_),
    .I1(_0475_),
    .S(_0109_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1323_ (.I0(_0202_),
    .I1(_0476_),
    .S(_0235_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1324_ (.A1(_0197_),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1325_ (.I0(_0230_),
    .I1(_0240_),
    .S(_0330_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1326_ (.A1(_0197_),
    .A2(_0479_),
    .B(_0074_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1327_ (.I0(_0091_),
    .I1(_0051_),
    .S(_0805_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1328_ (.I0(_0458_),
    .I1(_0481_),
    .S(_0127_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1329_ (.A1(_0122_),
    .A2(_0248_),
    .B1(_0482_),
    .B2(_0223_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1330_ (.A1(_0152_),
    .A2(_0384_),
    .B(_0209_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1331_ (.A1(_0152_),
    .A2(_0483_),
    .B1(_0484_),
    .B2(_0279_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1332_ (.A1(_0246_),
    .A2(_0272_),
    .B(_0485_),
    .C(_0215_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1333_ (.A1(_0473_),
    .A2(_0478_),
    .B1(_0480_),
    .B2(_0486_),
    .ZN(net49));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1334_ (.A1(_0040_),
    .A2(_0279_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1335_ (.A1(_0487_),
    .A2(_0438_),
    .A3(_0439_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1336_ (.I0(net23),
    .I1(_0018_),
    .S(_0047_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1337_ (.I0(_0022_),
    .I1(_0489_),
    .S(_0175_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1338_ (.I0(_0005_),
    .I1(_0126_),
    .S(_0174_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1339_ (.I0(_0490_),
    .I1(_0491_),
    .S(_0208_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1340_ (.I0(_0019_),
    .I1(_0006_),
    .S(_0805_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1341_ (.I0(_0017_),
    .I1(_0493_),
    .S(_0175_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1342_ (.I0(_0295_),
    .I1(_0494_),
    .S(_0121_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1343_ (.I0(_0492_),
    .I1(_0495_),
    .S(_0152_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1344_ (.A1(_0038_),
    .A2(_0307_),
    .B1(_0496_),
    .B2(_0252_),
    .C(_0195_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1345_ (.I0(_0003_),
    .I1(_0102_),
    .I2(_0004_),
    .I3(_0098_),
    .S0(_0086_),
    .S1(_0087_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1346_ (.I0(_0323_),
    .I1(_0498_),
    .S(_0094_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1347_ (.I0(_0014_),
    .I1(_0019_),
    .I2(_0015_),
    .I3(_0006_),
    .S0(_0100_),
    .S1(_0105_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1348_ (.I0(net12),
    .I1(net23),
    .I2(_0021_),
    .I3(_0018_),
    .S0(_0107_),
    .S1(_0105_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1349_ (.I0(_0500_),
    .I1(_0501_),
    .S(_0109_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1350_ (.I0(_0499_),
    .I1(_0502_),
    .S(_0111_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1351_ (.I0(_0453_),
    .I1(_0503_),
    .S(_0114_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1352_ (.A1(_0072_),
    .A2(_0307_),
    .B(_0504_),
    .C(_0266_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1353_ (.A1(_0488_),
    .A2(_0497_),
    .B(_0505_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1354_ (.A1(_0044_),
    .A2(_0167_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1355_ (.A1(_0810_),
    .A2(_0063_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1356_ (.A1(_0133_),
    .A2(_0721_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1357_ (.A1(_0508_),
    .A2(_0340_),
    .B(_0234_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1358_ (.A1(_0507_),
    .A2(_0509_),
    .B(_0050_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1359_ (.A1(_0506_),
    .A2(_0510_),
    .B(_0162_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1360_ (.I(_0048_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1361_ (.A1(_0193_),
    .A2(_0285_),
    .B(_0057_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _1362_ (.A1(_0162_),
    .A2(_0512_),
    .A3(_0358_),
    .B(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1363_ (.I0(_0253_),
    .I1(_0258_),
    .S(_0011_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1364_ (.A1(_0034_),
    .A2(_0041_),
    .A3(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1365_ (.A1(_0732_),
    .A2(_0752_),
    .B(_0208_),
    .C(_0792_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1366_ (.I0(_0082_),
    .I1(_0090_),
    .S(_0023_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1367_ (.I0(_0481_),
    .I1(_0518_),
    .S(_0000_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1368_ (.I0(_0409_),
    .I1(_0519_),
    .S(_0011_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1369_ (.A1(_0517_),
    .A2(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1370_ (.A1(_0800_),
    .A2(_0208_),
    .A3(_0262_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1371_ (.A1(net38),
    .A2(_0516_),
    .A3(_0521_),
    .A4(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _1372_ (.A1(_0511_),
    .A2(_0514_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1373_ (.I0(_0082_),
    .I1(_0090_),
    .S(_0139_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1374_ (.I0(_0474_),
    .I1(_0525_),
    .S(_0127_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1375_ (.I0(_0421_),
    .I1(_0526_),
    .S(_0228_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1376_ (.I0(_0289_),
    .I1(_0527_),
    .S(_0185_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1377_ (.A1(_0229_),
    .A2(_0080_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1378_ (.I0(_0268_),
    .I1(_0529_),
    .S(_0330_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _1379_ (.A1(_0511_),
    .A2(_0514_),
    .A3(_0528_),
    .B1(_0530_),
    .B2(_0523_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1380_ (.A1(_0337_),
    .A2(_0524_),
    .B(_0531_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1381_ (.I0(_0083_),
    .I1(_0091_),
    .S(_0047_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1382_ (.I0(_0518_),
    .I1(_0532_),
    .S(_0001_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1383_ (.I0(_0408_),
    .I1(_0431_),
    .S(_0001_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1384_ (.I0(_0533_),
    .I1(_0534_),
    .S(_0151_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1385_ (.I0(_0318_),
    .I1(_0535_),
    .S(_0223_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1386_ (.A1(_0215_),
    .A2(_0035_),
    .A3(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1387_ (.I0(_0333_),
    .I1(_0327_),
    .S(_0330_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1388_ (.A1(_0210_),
    .A2(_0320_),
    .B1(_0538_),
    .B2(_0132_),
    .C(_0266_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1389_ (.A1(_0012_),
    .A2(_0299_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1390_ (.I0(_0294_),
    .I1(_0540_),
    .S(_0209_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1391_ (.I0(_0083_),
    .I1(_0091_),
    .S(_0139_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1392_ (.I0(_0525_),
    .I1(_0542_),
    .S(_0662_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1393_ (.I0(_0445_),
    .I1(_0543_),
    .S(_0094_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1394_ (.I0(_0313_),
    .I1(_0544_),
    .S(_0234_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1395_ (.A1(_0185_),
    .A2(_0309_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1396_ (.I0(_0545_),
    .I1(_0546_),
    .S(_0328_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1397_ (.A1(_0802_),
    .A2(_0541_),
    .B(_0547_),
    .C(_0059_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1398_ (.A1(_0537_),
    .A2(_0539_),
    .B(_0548_),
    .ZN(net52));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _1399_ (.I(_0369_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1400_ (.A1(_0027_),
    .A2(_0118_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1401_ (.I0(_0345_),
    .I1(_0550_),
    .S(_0208_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1402_ (.A1(_0193_),
    .A2(_0549_),
    .B1(_0551_),
    .B2(_0802_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1403_ (.I0(_0166_),
    .I1(_0348_),
    .S(_0012_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1404_ (.I0(_0352_),
    .I1(_0354_),
    .S(_0150_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1405_ (.I0(_0084_),
    .I1(_0082_),
    .S(_0805_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1406_ (.I0(_0431_),
    .I1(_0458_),
    .I2(_0532_),
    .I3(_0555_),
    .S0(_0672_),
    .S1(_0027_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1407_ (.I0(_0554_),
    .I1(_0556_),
    .S(_0121_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1408_ (.A1(_0122_),
    .A2(_0553_),
    .B1(_0557_),
    .B2(_0223_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1409_ (.A1(_0266_),
    .A2(_0792_),
    .A3(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1410_ (.A1(_0254_),
    .A2(_0117_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1411_ (.I0(_0364_),
    .I1(_0560_),
    .S(_0330_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1412_ (.I0(_0084_),
    .I1(net13),
    .S(_0139_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1413_ (.I0(_0542_),
    .I1(_0562_),
    .S(_0127_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1414_ (.I0(_0466_),
    .I1(_0563_),
    .S(_0228_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1415_ (.I0(_0371_),
    .I1(_0564_),
    .S(_0234_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1416_ (.I0(_0561_),
    .I1(_0565_),
    .S(_0073_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1417_ (.A1(_0197_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _1418_ (.A1(_0059_),
    .A2(_0552_),
    .B(_0559_),
    .C(_0567_),
    .ZN(net53));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1419_ (.I0(net16),
    .I1(net14),
    .S(_0139_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1420_ (.I0(_0562_),
    .I1(_0568_),
    .S(_0662_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1421_ (.I0(_0475_),
    .I1(_0569_),
    .S(_0094_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1422_ (.I0(_0395_),
    .I1(_0570_),
    .S(_0235_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1423_ (.A1(_0330_),
    .A2(_0229_),
    .A3(net25),
    .A4(_0068_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1424_ (.A1(_0235_),
    .A2(_0398_),
    .B(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1425_ (.A1(_0073_),
    .A2(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1426_ (.A1(_0402_),
    .A2(_0571_),
    .B(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1427_ (.I0(_0085_),
    .I1(_0083_),
    .S(_0023_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1428_ (.I0(_0555_),
    .I1(_0576_),
    .S(_0127_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1429_ (.I0(_0384_),
    .I1(_0577_),
    .S(_0033_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1430_ (.I0(_0245_),
    .I1(_0482_),
    .S(_0033_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1431_ (.I0(_0578_),
    .I1(_0579_),
    .S(_0151_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1432_ (.A1(_0034_),
    .A2(_0381_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1433_ (.I0(_0580_),
    .I1(_0581_),
    .S(_0279_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1434_ (.A1(_0215_),
    .A2(_0582_),
    .B(_0074_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1435_ (.A1(_0027_),
    .A2(_0216_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1436_ (.I0(_0375_),
    .I1(_0584_),
    .S(_0208_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1437_ (.A1(_0193_),
    .A2(_0391_),
    .B1(_0585_),
    .B2(_0801_),
    .C(_0058_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _1438_ (.A1(_0337_),
    .A2(_0575_),
    .B1(_0583_),
    .B2(_0586_),
    .ZN(net54));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1439_ (.I0(_0403_),
    .I1(_0405_),
    .S(_0175_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1440_ (.A1(_0027_),
    .A2(_0253_),
    .A3(_0255_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1441_ (.A1(_0035_),
    .A2(_0587_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1442_ (.A1(_0487_),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1443_ (.A1(_0113_),
    .A2(_0096_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1444_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1445_ (.I0(_0153_),
    .I1(_0084_),
    .S(_0016_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1446_ (.I0(_0576_),
    .I1(_0593_),
    .S(_0672_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1447_ (.I0(_0409_),
    .I1(_0594_),
    .S(_0121_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1448_ (.I0(_0411_),
    .I1(_0519_),
    .S(_0121_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1449_ (.I0(_0595_),
    .I1(_0596_),
    .S(_0152_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1450_ (.A1(_0081_),
    .A2(_0592_),
    .B1(_0252_),
    .B2(_0597_),
    .C(_0266_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1451_ (.I(_0517_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1452_ (.A1(_0056_),
    .A2(_0254_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1453_ (.I0(_0419_),
    .I1(_0600_),
    .S(_0062_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1454_ (.I0(_0153_),
    .I1(net15),
    .S(_0139_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1455_ (.I0(_0568_),
    .I1(_0602_),
    .S(_0662_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1456_ (.I0(_0526_),
    .I1(_0603_),
    .S(_0109_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1457_ (.I0(_0422_),
    .I1(_0604_),
    .S(_0111_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1458_ (.I0(_0601_),
    .I1(_0605_),
    .S(_0114_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1459_ (.A1(_0049_),
    .A2(_0599_),
    .B(_0606_),
    .C(_0059_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1460_ (.A1(_0590_),
    .A2(_0598_),
    .B(_0607_),
    .ZN(net55));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1461_ (.A1(_0592_),
    .A2(_0451_),
    .B(_0402_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1462_ (.I0(_0045_),
    .I1(_0085_),
    .S(_0024_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1463_ (.I0(_0593_),
    .I1(_0609_),
    .S(_0001_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1464_ (.I0(_0533_),
    .I1(_0610_),
    .S(_0012_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1465_ (.I0(_0433_),
    .I1(_0611_),
    .S(_0035_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1466_ (.A1(_0167_),
    .A2(_0316_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1467_ (.A1(_0035_),
    .A2(_0427_),
    .B(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1468_ (.A1(_0487_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1469_ (.A1(_0802_),
    .A2(_0612_),
    .B(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1470_ (.A1(_0330_),
    .A2(_0254_),
    .A3(_0307_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1471_ (.A1(_0185_),
    .A2(_0443_),
    .B(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1472_ (.I0(_0045_),
    .I1(_0085_),
    .S(_0692_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1473_ (.I0(_0602_),
    .I1(_0619_),
    .S(_0672_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1474_ (.I0(_0312_),
    .I1(_0445_),
    .I2(_0543_),
    .I3(_0620_),
    .S0(_0203_),
    .S1(_0234_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1475_ (.A1(_0328_),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1476_ (.A1(_0337_),
    .A2(_0618_),
    .B(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1477_ (.A1(_0437_),
    .A2(_0599_),
    .B(_0623_),
    .C(_0195_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1478_ (.A1(_0608_),
    .A2(_0616_),
    .B(_0624_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1479_ (.I0(_0046_),
    .I1(_0153_),
    .S(_0016_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1480_ (.I0(_0532_),
    .I1(_0555_),
    .I2(_0609_),
    .I3(_0625_),
    .S0(_0808_),
    .S1(_0028_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1481_ (.I0(_0460_),
    .I1(_0626_),
    .S(_0035_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1482_ (.A1(_0802_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1483_ (.A1(_0487_),
    .A2(_0178_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1484_ (.A1(_0592_),
    .A2(_0191_),
    .B(_0629_),
    .C(_0074_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1485_ (.I0(_0046_),
    .I1(_0153_),
    .S(_0139_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1486_ (.I0(_0619_),
    .I1(_0631_),
    .S(_0127_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1487_ (.I0(_0563_),
    .I1(_0632_),
    .S(_0109_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1488_ (.I0(_0467_),
    .I1(_0633_),
    .S(_0111_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1489_ (.I0(_0148_),
    .I1(_0634_),
    .S(_0114_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1490_ (.A1(_0120_),
    .A2(_0599_),
    .B(_0635_),
    .C(_0195_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1491_ (.A1(_0628_),
    .A2(_0630_),
    .B(_0636_),
    .ZN(net57));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1492_ (.A1(_0592_),
    .A2(_0240_),
    .B1(_0250_),
    .B2(_0042_),
    .C(_0074_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1493_ (.I0(net20),
    .I1(_0045_),
    .S(_0016_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1494_ (.I0(_0625_),
    .I1(_0638_),
    .S(_0672_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1495_ (.I0(_0482_),
    .I1(_0639_),
    .S(_0121_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1496_ (.I0(_0578_),
    .I1(_0640_),
    .S(_0028_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1497_ (.A1(_0802_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1498_ (.I0(net20),
    .I1(_0045_),
    .S(_0692_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1499_ (.I0(_0631_),
    .I1(_0644_),
    .S(_0662_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1500_ (.I0(_0569_),
    .I1(_0645_),
    .S(_0109_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1501_ (.I0(_0476_),
    .I1(_0646_),
    .S(_0111_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1502_ (.I0(_0207_),
    .I1(_0647_),
    .S(_0114_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1503_ (.A1(_0218_),
    .A2(_0599_),
    .B(_0648_),
    .C(_0195_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1504_ (.A1(_0637_),
    .A2(_0643_),
    .B(_0649_),
    .ZN(net58));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1505_ (.A1(_0229_),
    .A2(_0592_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1506_ (.A1(_0042_),
    .A2(_0264_),
    .B1(_0650_),
    .B2(_0080_),
    .C(_0074_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1507_ (.I0(_0043_),
    .I1(_0046_),
    .S(_0024_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1508_ (.I0(_0638_),
    .I1(_0653_),
    .S(_0001_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1509_ (.I0(_0519_),
    .I1(_0654_),
    .S(_0034_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1510_ (.I0(_0595_),
    .I1(_0655_),
    .S(_0028_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1511_ (.A1(_0802_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1512_ (.I0(_0043_),
    .I1(_0046_),
    .S(_0692_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1513_ (.I0(_0644_),
    .I1(_0658_),
    .S(_0000_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1514_ (.I0(_0603_),
    .I1(_0659_),
    .S(_0228_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1515_ (.I0(_0527_),
    .I1(_0660_),
    .S(_0234_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1516_ (.I0(_0290_),
    .I1(_0661_),
    .S(_0132_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1517_ (.A1(_0071_),
    .A2(_0801_),
    .A3(_0044_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _1518_ (.A1(_0059_),
    .A2(_0663_),
    .A3(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1519_ (.A1(_0652_),
    .A2(_0657_),
    .B(_0665_),
    .ZN(net59));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1520_ (.I0(net22),
    .I1(net20),
    .S(_0024_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1521_ (.I0(_0593_),
    .I1(_0609_),
    .I2(_0653_),
    .I3(_0666_),
    .S0(_0808_),
    .S1(_0012_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1522_ (.I0(_0535_),
    .I1(_0667_),
    .S(_0035_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1523_ (.A1(_0042_),
    .A2(_0321_),
    .B1(_0668_),
    .B2(_0802_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1524_ (.A1(_0650_),
    .A2(_0326_),
    .B(_0402_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1525_ (.I0(net22),
    .I1(net20),
    .S(_0140_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1526_ (.I0(_0602_),
    .I1(_0619_),
    .I2(_0658_),
    .I3(_0671_),
    .S0(_0672_),
    .S1(_0228_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1527_ (.I0(_0544_),
    .I1(_0673_),
    .S(_0111_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1528_ (.I0(_0314_),
    .I1(_0674_),
    .S(_0114_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1529_ (.A1(_0599_),
    .A2(_0540_),
    .B(_0675_),
    .C(_0195_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1530_ (.A1(_0669_),
    .A2(_0670_),
    .B(_0676_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1531_ (.A1(_0133_),
    .A2(_0742_),
    .A3(_0146_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1532_ (.I0(_0021_),
    .I1(_0014_),
    .S(_0007_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1533_ (.I0(_0489_),
    .I1(_0678_),
    .S(_0174_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1534_ (.I0(_0128_),
    .I1(_0679_),
    .S(_0033_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1535_ (.I0(_0015_),
    .I1(net32),
    .S(_0804_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1536_ (.I0(_0493_),
    .I1(_0681_),
    .S(_0107_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1537_ (.I0(_0157_),
    .I1(_0682_),
    .S(_0033_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1538_ (.I0(_0680_),
    .I1(_0683_),
    .S(_0151_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1539_ (.A1(_0042_),
    .A2(_0464_),
    .B1(_0684_),
    .B2(_0801_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1540_ (.A1(_0402_),
    .A2(_0677_),
    .A3(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1541_ (.I0(_0019_),
    .I1(_0015_),
    .I2(_0006_),
    .I3(_0003_),
    .S0(_0067_),
    .S1(_0140_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1542_ (.I0(net23),
    .I1(_0021_),
    .I2(_0018_),
    .I3(_0014_),
    .S0(_0067_),
    .S1(_0140_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1543_ (.I0(_0687_),
    .I1(_0688_),
    .S(_0093_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1544_ (.I0(_0184_),
    .I1(_0689_),
    .S(_0096_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1545_ (.I0(_0455_),
    .I1(_0690_),
    .S(_0114_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1546_ (.A1(_0071_),
    .A2(_0800_),
    .A3(_0166_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1547_ (.A1(_0073_),
    .A2(_0691_),
    .A3(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1548_ (.A1(_0686_),
    .A2(_0694_),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1549_ (.A1(_0354_),
    .A2(_0358_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1550_ (.A1(_0487_),
    .A2(_0350_),
    .A3(_0353_),
    .A4(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1551_ (.I0(net24),
    .I1(_0043_),
    .S(_0024_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1552_ (.I0(_0609_),
    .I1(_0625_),
    .I2(_0666_),
    .I3(_0697_),
    .S0(_0808_),
    .S1(_0012_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1553_ (.I0(_0556_),
    .I1(_0698_),
    .S(_0177_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1554_ (.A1(_0038_),
    .A2(_0117_),
    .B1(_0699_),
    .B2(_0252_),
    .C(_0266_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1555_ (.A1(_0328_),
    .A2(_0373_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1556_ (.I0(net24),
    .I1(_0043_),
    .S(_0140_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1557_ (.I0(_0619_),
    .I1(_0631_),
    .I2(_0671_),
    .I3(_0702_),
    .S0(_0001_),
    .S1(_0203_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1558_ (.I0(_0564_),
    .I1(_0703_),
    .S(_0234_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1559_ (.A1(_0328_),
    .A2(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1560_ (.A1(_0072_),
    .A2(_0117_),
    .B1(_0701_),
    .B2(_0705_),
    .C(_0195_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1561_ (.A1(_0696_),
    .A2(_0700_),
    .B(_0706_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1562_ (.A1(_0245_),
    .A2(_0358_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1563_ (.A1(_0487_),
    .A2(_0382_),
    .A3(_0385_),
    .A4(_0707_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1564_ (.I0(net25),
    .I1(net24),
    .I2(net22),
    .I3(_0043_),
    .S0(_0174_),
    .S1(_0024_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1565_ (.I0(_0577_),
    .I1(_0709_),
    .S(_0121_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1566_ (.I0(_0640_),
    .I1(_0710_),
    .S(_0028_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1567_ (.A1(_0038_),
    .A2(_0387_),
    .B1(_0712_),
    .B2(_0252_),
    .C(_0266_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1568_ (.I0(net25),
    .I1(net24),
    .I2(net22),
    .I3(_0043_),
    .S0(_0107_),
    .S1(_0105_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1569_ (.I0(_0645_),
    .I1(_0714_),
    .S(_0109_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1570_ (.I0(_0570_),
    .I1(_0715_),
    .S(_0111_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1571_ (.I0(_0396_),
    .I1(_0716_),
    .S(_0114_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1572_ (.A1(_0072_),
    .A2(_0387_),
    .B(_0717_),
    .C(_0195_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1573_ (.A1(_0708_),
    .A2(_0713_),
    .B(_0718_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1574_ (.I0(_0233_),
    .I1(_0240_),
    .S(_0328_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1575_ (.I0(_0015_),
    .I1(_0006_),
    .I2(_0003_),
    .I3(_0102_),
    .S0(_0107_),
    .S1(_0105_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1576_ (.I0(_0021_),
    .I1(_0018_),
    .I2(_0014_),
    .I3(_0019_),
    .S0(_0175_),
    .S1(_0105_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1577_ (.I0(_0720_),
    .I1(_0722_),
    .S(_0229_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1578_ (.A1(_0592_),
    .A2(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1579_ (.A1(_0193_),
    .A2(_0230_),
    .B1(_0719_),
    .B2(_0330_),
    .C(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1580_ (.A1(_0071_),
    .A2(_0801_),
    .A3(_0248_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1581_ (.A1(_0402_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1582_ (.I0(_0008_),
    .I1(_0681_),
    .S(_0037_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1583_ (.I0(_0020_),
    .I1(_0678_),
    .S(_0662_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1584_ (.I0(_0728_),
    .I1(_0729_),
    .S(_0011_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1585_ (.I0(_0222_),
    .I1(_0730_),
    .S(_0121_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1586_ (.I0(_0472_),
    .I1(_0731_),
    .S(_0223_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1587_ (.A1(_0205_),
    .A2(_0650_),
    .B1(_0733_),
    .B2(_0215_),
    .C(_0058_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1588_ (.A1(_0725_),
    .A2(_0727_),
    .B(_0734_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1589_ (.I0(_0103_),
    .I1(_0106_),
    .S(_0203_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1590_ (.I0(_0269_),
    .I1(_0735_),
    .S(_0185_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1591_ (.A1(_0132_),
    .A2(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1592_ (.A1(_0337_),
    .A2(_0530_),
    .B(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1593_ (.A1(_0515_),
    .A2(_0599_),
    .B(_0402_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1594_ (.A1(_0592_),
    .A2(_0285_),
    .B(_0059_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _1595_ (.A1(_0512_),
    .A2(_0358_),
    .B(_0506_),
    .C(_0510_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1596_ (.I0(_0017_),
    .I1(_0020_),
    .S(_0808_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _1597_ (.I0(_0052_),
    .I1(_0002_),
    .I2(_0009_),
    .I3(_0743_),
    .S0(_0028_),
    .S1(_0177_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1598_ (.A1(_0042_),
    .A2(_0741_),
    .B1(_0744_),
    .B2(_0252_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1599_ (.A1(_0738_),
    .A2(_0739_),
    .B1(_0740_),
    .B2(_0745_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1600_ (.I0(_0498_),
    .I1(_0500_),
    .S(_0203_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1601_ (.I0(_0324_),
    .I1(_0746_),
    .S(_0185_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1602_ (.A1(_0132_),
    .A2(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1603_ (.A1(_0337_),
    .A2(_0538_),
    .B(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1604_ (.A1(_0318_),
    .A2(_0599_),
    .B(_0074_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1605_ (.A1(_0592_),
    .A2(_0309_),
    .B(_0059_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1606_ (.I0(_0301_),
    .I1(_0491_),
    .S(_0033_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1607_ (.I0(_0495_),
    .I1(_0753_),
    .S(_0152_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1608_ (.A1(_0042_),
    .A2(_0541_),
    .B1(_0754_),
    .B2(_0252_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _1609_ (.A1(_0749_),
    .A2(_0750_),
    .B1(_0751_),
    .B2(_0755_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1610_ (.I0(_0183_),
    .I1(_0687_),
    .S(_0228_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1611_ (.I0(_0365_),
    .I1(_0756_),
    .S(_0234_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1612_ (.I0(_0561_),
    .I1(_0757_),
    .S(_0132_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1613_ (.A1(_0553_),
    .A2(_0599_),
    .B(_0758_),
    .C(_0402_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1614_ (.I0(_0129_),
    .I1(_0683_),
    .S(_0012_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1615_ (.I0(_0551_),
    .I1(_0760_),
    .S(_0223_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1616_ (.A1(_0592_),
    .A2(_0549_),
    .B1(_0761_),
    .B2(_0215_),
    .C(_0059_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1617_ (.A1(_0759_),
    .A2(_0763_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1618_ (.I0(_0221_),
    .I1(_0728_),
    .S(_0011_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1619_ (.I0(_0378_),
    .I1(_0764_),
    .S(_0034_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1620_ (.I0(_0585_),
    .I1(_0765_),
    .S(_0223_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1621_ (.A1(_0592_),
    .A2(_0391_),
    .B1(_0766_),
    .B2(_0215_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1622_ (.I0(_0232_),
    .I1(_0720_),
    .S(_0228_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1623_ (.I0(_0399_),
    .I1(_0768_),
    .S(_0234_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1624_ (.A1(_0328_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1625_ (.A1(_0328_),
    .A2(_0573_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _1626_ (.A1(_0381_),
    .A2(_0599_),
    .B(_0771_),
    .C(_0266_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _1627_ (.A1(_0402_),
    .A2(_0767_),
    .B(_0773_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1628_ (.I0(_0050_),
    .I1(_0002_),
    .S(_0034_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1629_ (.A1(_0028_),
    .A2(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1630_ (.I(_0052_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1631_ (.A1(_0064_),
    .A2(_0070_),
    .B(_0009_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1632_ (.A1(_0776_),
    .A2(_0167_),
    .B(_0777_),
    .C(_0162_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1633_ (.A1(_0177_),
    .A2(_0049_),
    .A3(_0042_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1634_ (.A1(_0058_),
    .A2(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1635_ (.A1(_0197_),
    .A2(_0601_),
    .B1(_0775_),
    .B2(_0778_),
    .C(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1636_ (.I0(_0095_),
    .I1(_0104_),
    .S(_0185_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1637_ (.A1(_0599_),
    .A2(_0587_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1638_ (.A1(_0800_),
    .A2(_0588_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _1639_ (.A1(_0073_),
    .A2(_0784_),
    .A3(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1640_ (.A1(_0081_),
    .A2(_0193_),
    .B1(_0783_),
    .B2(_0132_),
    .C(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _1641_ (.A1(_0781_),
    .A2(_0787_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1642_ (.I0(_0295_),
    .I1(_0292_),
    .S(_0208_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1643_ (.I0(_0753_),
    .I1(_0788_),
    .S(_0151_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1644_ (.A1(_0034_),
    .A2(_0041_),
    .A3(_0437_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _1645_ (.A1(_0801_),
    .A2(_0789_),
    .B(_0790_),
    .C(_0058_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1646_ (.A1(_0193_),
    .A2(_0451_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _1647_ (.A1(_0427_),
    .A2(_0517_),
    .B1(_0613_),
    .B2(_0800_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1648_ (.A1(_0058_),
    .A2(_0793_),
    .A3(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1649_ (.A1(_0791_),
    .A2(_0795_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1650_ (.A1(_0330_),
    .A2(_0452_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1651_ (.A1(_0235_),
    .A2(_0499_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1652_ (.A1(_0795_),
    .A2(_0797_),
    .A3(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _1653_ (.A1(_0618_),
    .A2(_0791_),
    .B1(_0796_),
    .B2(_0337_),
    .C(_0799_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _1654_ (.A(_0808_),
    .B(_0809_),
    .CO(_0810_),
    .S(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Right_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Right_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Right_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Right_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Right_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Right_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Right_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Right_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Right_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Right_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Right_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Right_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Right_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Right_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Right_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Right_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Right_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Right_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Right_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Right_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Right_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Right_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Right_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Right_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Right_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Right_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Right_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Right_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Right_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Right_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Right_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Right_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Right_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Right_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Right_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Right_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Right_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Right_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Right_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Right_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Right_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Right_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Right_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Right_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Right_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Right_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Right_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Right_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Right_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Right_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Right_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Right_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Right_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Right_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Right_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Right_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Right_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Right_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Right_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Right_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Right_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Right_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Right_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Right_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Right_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Right_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Right_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Right_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Right_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Right_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Right_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Right_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Right_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Right_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Right_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Right_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Right_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Right_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Right_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Right_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Right_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Right_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Right_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Right_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Right_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Right_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Right_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Right_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Right_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Right_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Right_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Right_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Right_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Right_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Right_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Right_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_342_Right_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_343_Right_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_344_Right_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_345_Right_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_346_Right_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_347_Right_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_348_Right_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_349_Right_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_350_Right_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_351_Right_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_352_Right_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_353_Right_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_354_Right_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_355_Right_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_356_Right_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_357_Right_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_358_Right_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_359_Right_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_360_Right_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_361_Right_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_362_Right_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_363_Right_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_364_Right_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_365_Right_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_366_Right_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_367_Right_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_368_Right_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_369_Right_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_370_Right_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_371_Right_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_372_Right_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_373_Right_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_374_Right_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_375_Right_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_376_Right_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_377_Right_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_378_Right_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_379_Right_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_380_Right_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_381_Right_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_382_Right_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_383_Right_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_384_Right_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_385_Right_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_386_Right_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_387_Right_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_388_Right_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_389_Right_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_390_Right_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_391_Right_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_392_Right_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_393_Right_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_394_Right_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_395_Right_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_396_Right_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_397_Right_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_398_Right_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_399_Right_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_400_Right_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_401_Right_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_402_Right_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_403_Right_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_404_Right_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_405_Right_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_406_Right_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_407_Right_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_408_Right_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_409_Right_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_410_Right_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_411_Right_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_412_Right_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_413_Right_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_414_Right_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_415_Right_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_416_Right_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_417_Right_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_418_Right_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_419_Right_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_420_Right_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_421_Right_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_422_Right_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_423_Right_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_424_Right_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_425_Right_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_426_Right_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_427_Right_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_428_Right_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_429_Right_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_430_Right_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_431_Right_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_432_Right_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_433_Right_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_434_Right_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_435_Right_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_436_Right_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_437_Right_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_438_Right_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_439_Right_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_440_Right_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_441_Right_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_442_Right_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_443_Right_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_444_Right_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_445_Right_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_446_Right_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_447_Right_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_448_Right_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_449_Right_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_450_Right_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_451_Right_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_452_Right_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_453_Right_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_454_Right_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_455_Right_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_456_Right_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_457_Right_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_458_Right_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_459_Right_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_460_Right_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_461_Right_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_462_Right_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_463_Right_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_464_Right_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_465_Right_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_466_Right_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_467_Right_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_468_Right_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_469_Right_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_470_Right_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_471_Right_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_472_Right_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_473_Right_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_474_Right_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_475_Right_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_476_Right_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_477_Right_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_478_Right_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_479_Right_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_480_Right_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_481_Right_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_482_Right_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_483_Right_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_484_Right_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_485_Right_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_486_Right_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_487_Right_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_488_Right_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_489_Right_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_490_Right_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_491_Right_491 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_492_Right_492 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_493_Right_493 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_494_Right_494 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_495_Right_495 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_496_Right_496 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_497_Right_497 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_498_Right_498 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_499_Right_499 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_500_Right_500 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_501_Right_501 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_502_Right_502 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_503_Right_503 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_504_Right_504 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_505_Right_505 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_506_Right_506 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_507 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_508 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_509 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_510 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_511 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_512 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_513 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_514 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_515 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_516 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_517 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_518 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_519 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_520 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_521 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_522 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_523 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_524 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_525 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_526 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_527 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_528 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_529 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_530 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_531 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_532 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_533 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_534 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_535 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_536 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_537 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_538 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_539 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_540 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_541 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_542 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_543 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_544 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_545 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_546 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_547 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_548 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_549 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_550 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_551 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_552 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_553 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_554 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_555 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_556 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_557 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_558 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_559 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_560 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_561 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_562 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_563 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_564 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_565 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_566 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_567 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_568 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_569 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_570 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_571 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_572 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_573 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_574 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_575 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_576 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_577 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_578 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_579 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_580 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_581 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_582 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_583 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_584 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_585 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_586 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_587 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_588 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_589 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_590 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_591 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_592 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_593 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_594 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_595 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_596 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_597 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_598 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_599 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_600 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_601 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_602 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_603 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_604 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_605 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_606 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_607 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_608 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_609 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_610 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_611 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_612 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_613 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_614 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_615 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_616 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_617 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_618 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_619 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_620 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_621 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_622 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_623 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_624 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_625 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_626 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_627 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_628 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_629 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_630 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_631 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_632 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_633 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_634 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_635 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_636 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_637 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_638 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_639 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_640 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_641 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_642 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_643 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_644 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_645 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_646 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_647 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_648 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_649 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_650 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_651 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_652 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_653 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_654 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_655 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_656 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_657 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_658 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_659 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_660 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_661 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_662 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_663 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_664 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_665 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_666 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_667 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_668 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_669 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_670 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_671 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_672 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_673 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_674 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_675 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_676 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_677 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_678 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_679 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_680 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_681 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_682 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_683 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_684 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_685 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_686 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_687 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_688 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_689 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_690 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_691 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_692 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_693 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_694 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_695 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_696 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_697 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_698 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_699 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_700 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_701 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_702 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_703 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_704 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_705 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_706 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_707 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_708 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_709 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_710 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_711 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_712 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_713 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_714 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_715 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_716 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_717 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_718 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_719 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_720 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_721 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_722 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_723 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_724 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_725 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_726 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_727 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_728 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_729 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_730 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_731 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_732 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_733 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_734 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_735 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_736 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_737 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_738 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_739 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_740 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_741 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_742 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_743 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_744 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_745 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_746 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_747 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_748 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_749 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_750 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_751 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_752 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Left_753 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Left_754 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Left_755 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Left_756 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Left_757 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Left_758 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Left_759 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Left_760 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Left_761 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Left_762 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Left_763 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Left_764 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Left_765 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Left_766 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Left_767 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Left_768 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Left_769 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Left_770 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Left_771 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Left_772 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Left_773 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Left_774 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Left_775 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Left_776 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Left_777 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Left_778 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Left_779 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Left_780 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Left_781 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Left_782 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Left_783 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Left_784 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Left_785 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Left_786 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Left_787 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Left_788 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Left_789 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Left_790 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Left_791 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Left_792 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Left_793 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Left_794 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Left_795 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Left_796 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Left_797 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Left_798 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Left_799 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Left_800 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Left_801 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Left_802 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Left_803 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Left_804 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Left_805 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Left_806 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Left_807 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Left_808 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Left_809 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Left_810 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Left_811 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Left_812 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Left_813 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Left_814 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Left_815 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Left_816 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Left_817 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Left_818 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Left_819 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Left_820 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Left_821 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Left_822 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Left_823 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Left_824 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Left_825 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Left_826 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Left_827 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Left_828 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Left_829 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Left_830 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Left_831 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Left_832 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Left_833 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Left_834 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Left_835 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Left_836 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Left_837 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Left_838 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Left_839 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Left_840 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Left_841 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Left_842 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Left_843 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Left_844 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Left_845 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Left_846 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Left_847 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Left_848 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_342_Left_849 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_343_Left_850 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_344_Left_851 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_345_Left_852 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_346_Left_853 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_347_Left_854 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_348_Left_855 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_349_Left_856 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_350_Left_857 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_351_Left_858 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_352_Left_859 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_353_Left_860 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_354_Left_861 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_355_Left_862 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_356_Left_863 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_357_Left_864 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_358_Left_865 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_359_Left_866 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_360_Left_867 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_361_Left_868 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_362_Left_869 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_363_Left_870 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_364_Left_871 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_365_Left_872 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_366_Left_873 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_367_Left_874 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_368_Left_875 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_369_Left_876 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_370_Left_877 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_371_Left_878 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_372_Left_879 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_373_Left_880 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_374_Left_881 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_375_Left_882 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_376_Left_883 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_377_Left_884 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_378_Left_885 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_379_Left_886 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_380_Left_887 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_381_Left_888 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_382_Left_889 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_383_Left_890 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_384_Left_891 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_385_Left_892 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_386_Left_893 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_387_Left_894 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_388_Left_895 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_389_Left_896 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_390_Left_897 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_391_Left_898 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_392_Left_899 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_393_Left_900 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_394_Left_901 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_395_Left_902 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_396_Left_903 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_397_Left_904 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_398_Left_905 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_399_Left_906 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_400_Left_907 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_401_Left_908 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_402_Left_909 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_403_Left_910 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_404_Left_911 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_405_Left_912 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_406_Left_913 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_407_Left_914 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_408_Left_915 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_409_Left_916 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_410_Left_917 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_411_Left_918 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_412_Left_919 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_413_Left_920 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_414_Left_921 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_415_Left_922 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_416_Left_923 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_417_Left_924 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_418_Left_925 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_419_Left_926 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_420_Left_927 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_421_Left_928 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_422_Left_929 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_423_Left_930 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_424_Left_931 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_425_Left_932 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_426_Left_933 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_427_Left_934 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_428_Left_935 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_429_Left_936 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_430_Left_937 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_431_Left_938 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_432_Left_939 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_433_Left_940 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_434_Left_941 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_435_Left_942 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_436_Left_943 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_437_Left_944 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_438_Left_945 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_439_Left_946 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_440_Left_947 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_441_Left_948 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_442_Left_949 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_443_Left_950 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_444_Left_951 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_445_Left_952 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_446_Left_953 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_447_Left_954 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_448_Left_955 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_449_Left_956 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_450_Left_957 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_451_Left_958 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_452_Left_959 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_453_Left_960 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_454_Left_961 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_455_Left_962 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_456_Left_963 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_457_Left_964 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_458_Left_965 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_459_Left_966 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_460_Left_967 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_461_Left_968 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_462_Left_969 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_463_Left_970 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_464_Left_971 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_465_Left_972 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_466_Left_973 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_467_Left_974 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_468_Left_975 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_469_Left_976 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_470_Left_977 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_471_Left_978 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_472_Left_979 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_473_Left_980 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_474_Left_981 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_475_Left_982 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_476_Left_983 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_477_Left_984 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_478_Left_985 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_479_Left_986 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_480_Left_987 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_481_Left_988 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_482_Left_989 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_483_Left_990 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_484_Left_991 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_485_Left_992 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_486_Left_993 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_487_Left_994 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_488_Left_995 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_489_Left_996 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_490_Left_997 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_491_Left_998 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_492_Left_999 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_493_Left_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_494_Left_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_495_Left_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_496_Left_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_497_Left_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_498_Left_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_499_Left_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_500_Left_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_501_Left_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_502_Left_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_503_Left_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_504_Left_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_505_Left_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_506_Left_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_2225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_2325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_2338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_2400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_2488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_2513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_2538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_2563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_2588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_2625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_2638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_2675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_2688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_2700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_2713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_2725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_2738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_2763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_2775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_2788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_2813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_2825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_2838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_2863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_2875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_2888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_2900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_2913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_2925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_2938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_2950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_2963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_2975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_2988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_2999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_3000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_3013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_3025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_3038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_3050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_3063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_3075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_3088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_3100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_3113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_3125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_3138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_3150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_3163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_3175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_3200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_3213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_3225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_3238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_3250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_3263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_3275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_3288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_3300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_3313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_3325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_3338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_3350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_3363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_3375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_3388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_3400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_3413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_3425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_3438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_3450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_3463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_3475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_3488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_3500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_3513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_3525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_3538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_3550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_3563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_3575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_3588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_3600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_3613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_3625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_3638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_3650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_3663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_3675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_3688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_3700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_3713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_3725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_3738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_3750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_3763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_3775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_3788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_3800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_3813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_3825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_3838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_3850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_3863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_3875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_3888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_3913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_3925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_3938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_3950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_3963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_3975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_3988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_3999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_4000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_4013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_4025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_4038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_4050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_4063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_4075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_4088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_4100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_4113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_4125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_4138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_4150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_4163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_4175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_4188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_4200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_4213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_4225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_4250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_4263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_4275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_4300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_4313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_4325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_4350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_4363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_4375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_4388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_4400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_4413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_4425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_4438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_4450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_4463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_4475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_4488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_4500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_4513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_4525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_4538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_4550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_4563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_4575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_4588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_4600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_4613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_4625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_4638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_4650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_4663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_4675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_4688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_4700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_4713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_4725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_4738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_4750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_4763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_4775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_4788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_4800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_4813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_4825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_4838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_4850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_4863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_4875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_4888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_4900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_4913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_4925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_4938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_4950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_4963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_4975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_4988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_4999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_5000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_5013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_5025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_5038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_5050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_5063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_5075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_5088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_5100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_5113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_5125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_5138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_5150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_5163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_5175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_5188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_5200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_5213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_5225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_5238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_5250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_5263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_5275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_5288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_5300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_342_5313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_343_5325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_344_5338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_345_5350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_346_5363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_347_5375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_348_5388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_349_5400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_350_5413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_351_5425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_352_5438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_353_5450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_354_5463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_355_5475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_356_5488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_357_5500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_358_5513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_359_5525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_360_5538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_361_5550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_362_5563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_363_5575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_364_5588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_365_5600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_366_5613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_367_5625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_368_5638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_369_5650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_370_5663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_371_5675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_372_5688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_373_5700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_374_5713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_375_5725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_376_5738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_377_5750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_378_5763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_379_5775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_380_5788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_381_5800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_382_5813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_383_5825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_384_5838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_385_5850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_386_5863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_387_5875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_388_5888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_389_5900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_390_5913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_391_5925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_392_5938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_393_5950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_394_5963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_395_5975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_396_5988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_5999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_397_6000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_398_6013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_399_6025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_400_6038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_401_6050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_402_6063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_403_6075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_404_6088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_405_6100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_406_6113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_407_6125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_408_6138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_409_6150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_410_6163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_411_6175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_412_6188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_413_6200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_414_6213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_415_6225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_416_6238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_417_6250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_418_6263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_419_6275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_420_6288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_421_6300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_422_6313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_423_6325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_424_6338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_425_6350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_426_6363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_427_6375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_428_6388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_429_6400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_430_6413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_431_6425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_432_6438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_433_6450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_434_6463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_435_6475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_436_6488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_437_6500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_438_6513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_439_6525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_440_6538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_441_6550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_442_6563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_443_6575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_444_6588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_445_6600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_446_6613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_447_6625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_448_6638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_449_6650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_450_6663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_451_6675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_452_6688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_453_6700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_454_6713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_455_6725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_456_6738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_457_6750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_458_6763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_459_6775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_460_6788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_461_6800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_462_6813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_463_6825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_464_6838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_465_6850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_466_6863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_467_6875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_468_6888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_469_6900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_470_6913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_471_6925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_472_6938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_473_6950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_474_6963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_475_6975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_476_6988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_6999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_477_7000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_478_7013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_479_7025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_480_7038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_481_7050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_482_7063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_483_7075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_484_7088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_485_7100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_486_7113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_487_7125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_488_7138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_489_7150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_490_7163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_491_7175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_492_7188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_493_7200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_494_7213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_495_7225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_496_7238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_497_7250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_498_7263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_499_7275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_500_7288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_501_7300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_502_7313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_503_7325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_504_7338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_505_7350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_506_7375 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input1 (.I(data_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input2 (.I(data_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input3 (.I(data_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input4 (.I(data_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input5 (.I(data_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input6 (.I(data_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input7 (.I(data_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input8 (.I(data_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input9 (.I(data_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input10 (.I(data_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input11 (.I(data_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input12 (.I(data_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input13 (.I(data_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input14 (.I(data_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input15 (.I(data_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input16 (.I(data_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input17 (.I(data_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input18 (.I(data_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input19 (.I(data_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input20 (.I(data_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input21 (.I(data_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input22 (.I(data_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input23 (.I(data_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input24 (.I(data_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input25 (.I(data_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input26 (.I(data_in[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input27 (.I(data_in[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input28 (.I(data_in[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input29 (.I(data_in[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input30 (.I(data_in[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input31 (.I(data_in[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input32 (.I(data_in[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input33 (.I(rotate),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input34 (.I(shift_amount[1]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input35 (.I(shift_amount[2]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input36 (.I(shift_amount[3]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 input37 (.I(shift_amount[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input38 (.I(shift_direction),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net39),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net40),
    .Z(data_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net41),
    .Z(data_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net42),
    .Z(data_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net43),
    .Z(data_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net44),
    .Z(data_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net45),
    .Z(data_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net46),
    .Z(data_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net47),
    .Z(data_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net48),
    .Z(data_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net49),
    .Z(data_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net50),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net51),
    .Z(data_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net52),
    .Z(data_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net53),
    .Z(data_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net54),
    .Z(data_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net55),
    .Z(data_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net56),
    .Z(data_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net57),
    .Z(data_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net58),
    .Z(data_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net59),
    .Z(data_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net60),
    .Z(data_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net61),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net62),
    .Z(data_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net63),
    .Z(data_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net64),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net65),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(data_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(data_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net37));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net37));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net37));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_4078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_4256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_4434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_2492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_4506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_4508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_4547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_4563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_2660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_2649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_2259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_2361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_235_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_235_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_236_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_236_2412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_236_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_237_2839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_237_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_238_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_2647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_2422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_239_2467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_239_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_240_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_241_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_241_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_242_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_243_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_243_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_244_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_245_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_245_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_246_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_246_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_2666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_246_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_246_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_246_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_246_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_246_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_246_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_247_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_2274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_247_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_247_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_247_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_247_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_247_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_247_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_2230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_248_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_2648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_248_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_248_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_248_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_248_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_248_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_248_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_2539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_2811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_249_2843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_249_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_249_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_249_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_249_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_249_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_249_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_250_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_250_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_250_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_250_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_250_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_250_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_250_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_251_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_251_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_251_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_251_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_2809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_251_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_251_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_251_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_251_4518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_251_4533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_251_4565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_252_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_252_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_252_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_252_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_252_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_252_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_252_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_253_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_253_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_253_2517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_2796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_253_2828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_253_2844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_253_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_253_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_253_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_253_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_253_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_254_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_2429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_254_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_254_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_254_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_254_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_254_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_254_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_255_2440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_255_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_255_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_255_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_255_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_255_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_255_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_256_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_256_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_2428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_256_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_256_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_256_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_256_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_256_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_256_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_256_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_2425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_2817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_2833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_257_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_257_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_257_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_257_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_257_4543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_257_4559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_257_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_2300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_2409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_258_2519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_2645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_2661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_258_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_258_4484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_258_4500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_258_4508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_258_4535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_258_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_259_2424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_2809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_259_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_259_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_259_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_259_4498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_259_4514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_259_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_260_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_260_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_260_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_260_2482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_260_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_260_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_260_4520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_260_4547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_260_4563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_260_4567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_261_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_2518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_2807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_261_2839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_261_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_261_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_261_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_261_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_261_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_2236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_2643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_262_2659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_262_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_262_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_262_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_262_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_262_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_262_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_263_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_263_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_263_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_263_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_263_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_263_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_263_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_263_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_2359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_264_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_264_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_264_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_264_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_264_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_264_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_264_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_265_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_265_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_265_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_2431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_265_2464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_265_2480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_2488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_265_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_265_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_265_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_265_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_265_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_266_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_2650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_2666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_266_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_266_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_266_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_266_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_266_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_266_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_2303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_267_2433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_267_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_2457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_267_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_267_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_267_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_267_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_267_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_2286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_2495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_268_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_268_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_268_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_268_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_268_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_268_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_268_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_2351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_269_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_269_2481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_269_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_269_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_269_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_269_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_269_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_2505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_2509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_2646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_270_2662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_270_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_270_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_270_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_270_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_270_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_270_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_271_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_271_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_271_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_2506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_2843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_271_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_271_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_271_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_271_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_271_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_272_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_272_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_2640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_272_2656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_272_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_272_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_272_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_272_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_272_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_272_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_2294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_273_2475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_2805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_273_2837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_273_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_273_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_273_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_273_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_273_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_2260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_2340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_2456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_2641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_274_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_2665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_274_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_274_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_274_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_274_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_274_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_274_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_275_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_275_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_275_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_2253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_275_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_275_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_275_2384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_275_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_275_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_275_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_275_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_275_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_2196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_2250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_2284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_2292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_2419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_276_2435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_276_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_276_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_276_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_276_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_276_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_276_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_2267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_2785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_277_2817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_277_2833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_2841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_2845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_2847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_277_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_277_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_277_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_277_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_277_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_278_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_2208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_2227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_2248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_278_2396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_2664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_278_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_278_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_278_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_278_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_278_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_278_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_2252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_2256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_279_2272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_2304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_279_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_2399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_279_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_279_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_279_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_279_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_279_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_279_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_280_2299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_2307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_280_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_2401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_2417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_2653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_280_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_280_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_280_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_280_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_280_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_280_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_281_2283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_2360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_281_2462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_281_2478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_281_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_281_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_281_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_281_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_281_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_2354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_282_2402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_2651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_282_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_282_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_282_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_282_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_282_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_282_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_283_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_2329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_2335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_283_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_283_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_283_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_283_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_283_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_2341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_284_2347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_284_2363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_2639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_284_2655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_2663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_284_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_284_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_284_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_284_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_284_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_284_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_284_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_2308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_2324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_285_2339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_285_2355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_285_2484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_285_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_285_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_285_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_285_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_285_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_286_2661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_286_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_286_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_286_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_286_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_286_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_286_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_287_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_287_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_287_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_287_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_287_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_288_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_288_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_288_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_288_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_288_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_288_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_289_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_289_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_289_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_289_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_289_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_290_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_290_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_290_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_290_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_290_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_290_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_291_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_291_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_291_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_291_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_291_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_292_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_292_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_292_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_292_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_292_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_292_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_293_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_293_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_293_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_293_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_293_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_294_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_294_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_294_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_294_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_294_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_294_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_295_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_295_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_295_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_295_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_295_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_296_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_296_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_296_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_296_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_296_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_296_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_297_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_297_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_297_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_297_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_297_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_298_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_298_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_298_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_298_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_298_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_298_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_299_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_299_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_299_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_299_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_299_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_300_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_300_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_300_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_300_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_300_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_300_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_301_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_301_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_301_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_301_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_301_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_302_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_302_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_302_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_302_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_302_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_302_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_303_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_303_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_303_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_303_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_303_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_304_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_304_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_304_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_304_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_304_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_304_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_305_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_305_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_305_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_305_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_305_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_306_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_306_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_306_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_306_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_306_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_306_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_307_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_307_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_307_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_307_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_307_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_308_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_308_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_308_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_308_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_308_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_308_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_309_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_309_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_309_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_309_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_309_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_310_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_310_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_310_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_310_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_310_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_310_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_310_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_311_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_311_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_311_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_311_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_311_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_312_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_312_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_312_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_312_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_312_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_312_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_312_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_313_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_313_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_313_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_313_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_313_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_314_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_314_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_314_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_314_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_314_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_314_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_314_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_315_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_315_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_315_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_315_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_315_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_316_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_316_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_316_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_316_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_316_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_316_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_316_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_317_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_317_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_317_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_317_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_317_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_318_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_318_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_318_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_318_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_318_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_318_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_318_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_319_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_319_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_319_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_319_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_319_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_320_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_320_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_320_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_320_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_320_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_320_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_320_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_321_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_321_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_321_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_321_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_321_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_322_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_322_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_322_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_322_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_322_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_322_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_322_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_323_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_323_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_323_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_323_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_323_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_324_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_324_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_324_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_324_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_324_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_324_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_324_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_325_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_325_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_325_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_325_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_325_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_326_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_326_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_326_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_326_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_326_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_326_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_326_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_327_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_327_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_327_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_327_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_327_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_328_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_328_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_328_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_328_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_328_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_328_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_328_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_329_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_329_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_329_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_329_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_329_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_330_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_330_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_330_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_330_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_330_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_330_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_330_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_331_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_331_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_331_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_331_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_331_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_332_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_332_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_332_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_332_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_332_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_332_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_332_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_333_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_333_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_333_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_333_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_333_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_334_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_334_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_334_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_334_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_334_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_334_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_334_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_335_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_335_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_335_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_335_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_335_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_336_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_336_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_336_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_336_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_336_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_336_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_336_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_337_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_337_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_337_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_337_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_337_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_338_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_338_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_338_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_338_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_338_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_338_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_338_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_339_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_339_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_339_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_339_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_339_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_340_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_340_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_340_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_340_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_340_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_340_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_340_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_341_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_341_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_341_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_341_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_341_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_342_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_342_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_342_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_342_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_342_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_342_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_342_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_343_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_343_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_343_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_343_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_343_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_344_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_344_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_344_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_344_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_344_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_344_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_344_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_345_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_345_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_345_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_345_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_345_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_346_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_346_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_346_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_346_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_346_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_346_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_346_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_347_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_347_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_347_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_347_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_347_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_348_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_348_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_348_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_348_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_348_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_348_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_348_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_349_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_349_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_349_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_349_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_349_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_350_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_350_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_350_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_350_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_350_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_350_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_350_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_351_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_351_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_351_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_351_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_351_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_352_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_352_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_352_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_352_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_352_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_352_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_352_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_353_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_353_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_353_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_353_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_353_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_354_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_354_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_354_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_354_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_354_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_354_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_354_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_355_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_355_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_355_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_355_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_355_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_356_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_356_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_356_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_356_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_356_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_356_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_356_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_357_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_357_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_357_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_357_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_357_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_358_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_358_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_358_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_358_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_358_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_358_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_358_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_359_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_359_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_359_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_359_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_359_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_360_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_360_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_360_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_360_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_360_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_360_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_360_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_361_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_361_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_361_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_361_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_361_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_362_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_362_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_362_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_362_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_362_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_362_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_362_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_363_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_363_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_363_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_363_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_363_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_364_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_364_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_364_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_364_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_364_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_364_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_364_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_365_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_365_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_365_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_365_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_365_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_366_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_366_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_366_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_366_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_366_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_366_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_366_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_367_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_367_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_367_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_367_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_367_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_368_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_368_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_368_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_368_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_368_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_368_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_368_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_369_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_369_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_369_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_369_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_369_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_370_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_370_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_370_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_370_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_370_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_370_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_370_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_371_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_371_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_371_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_371_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_371_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_372_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_372_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_372_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_372_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_372_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_372_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_372_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_373_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_373_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_373_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_373_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_373_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_374_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_374_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_374_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_374_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_374_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_374_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_374_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_375_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_375_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_375_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_375_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_375_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_376_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_376_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_376_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_376_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_376_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_376_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_376_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_377_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_377_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_377_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_377_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_377_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_378_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_378_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_378_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_378_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_378_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_378_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_378_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_379_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_379_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_379_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_379_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_379_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_380_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_380_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_380_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_380_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_380_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_380_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_380_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_381_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_381_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_381_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_381_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_381_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_382_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_382_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_382_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_382_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_382_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_382_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_382_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_383_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_383_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_383_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_383_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_383_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_384_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_384_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_384_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_384_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_384_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_384_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_384_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_385_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_385_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_385_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_385_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_385_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_386_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_386_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_386_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_386_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_386_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_386_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_386_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_387_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_387_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_387_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_387_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_387_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_388_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_388_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_388_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_388_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_388_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_388_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_388_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_389_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_389_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_389_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_389_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_389_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_390_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_390_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_390_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_390_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_390_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_390_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_390_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_391_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_391_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_391_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_391_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_391_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_392_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_392_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_392_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_392_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_392_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_392_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_392_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_393_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_393_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_393_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_393_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_393_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_394_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_394_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_394_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_394_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_394_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_394_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_394_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_395_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_395_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_395_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_395_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_395_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_396_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_396_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_396_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_396_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_396_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_396_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_396_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_397_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_397_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_397_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_397_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_397_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_398_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_398_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_398_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_398_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_398_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_398_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_398_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_399_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_399_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_399_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_399_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_399_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_400_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_400_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_400_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_400_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_400_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_400_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_400_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_401_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_401_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_401_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_401_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_401_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_402_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_402_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_402_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_402_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_402_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_402_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_402_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_403_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_403_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_403_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_403_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_403_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_404_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_404_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_404_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_404_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_404_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_404_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_404_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_405_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_405_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_405_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_405_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_405_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_406_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_406_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_406_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_406_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_406_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_406_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_406_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_407_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_407_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_407_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_407_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_407_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_408_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_408_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_408_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_408_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_408_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_408_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_408_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_409_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_409_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_409_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_409_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_409_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_410_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_410_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_410_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_410_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_410_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_410_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_410_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_411_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_411_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_411_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_411_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_411_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_412_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_412_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_412_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_412_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_412_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_412_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_412_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_413_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_413_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_413_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_413_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_413_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_414_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_414_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_414_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_414_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_414_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_414_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_414_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_415_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_415_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_415_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_415_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_415_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_416_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_416_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_416_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_416_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_416_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_416_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_416_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_417_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_417_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_417_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_417_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_417_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_418_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_418_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_418_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_418_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_418_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_418_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_418_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_419_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_419_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_419_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_419_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_419_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_420_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_420_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_420_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_420_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_420_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_420_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_420_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_421_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_421_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_421_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_421_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_421_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_422_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_422_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_422_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_422_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_422_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_422_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_422_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_423_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_423_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_423_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_423_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_423_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_424_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_424_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_424_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_424_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_424_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_424_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_424_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_425_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_425_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_425_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_425_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_425_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_426_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_426_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_426_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_426_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_426_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_426_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_426_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_427_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_427_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_427_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_427_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_427_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_428_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_428_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_428_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_428_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_428_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_428_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_428_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_429_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_429_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_429_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_429_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_429_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_430_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_430_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_430_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_430_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_430_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_430_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_430_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_431_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_431_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_431_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_431_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_431_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_432_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_432_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_432_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_432_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_432_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_432_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_432_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_433_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_433_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_433_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_433_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_433_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_434_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_434_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_434_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_434_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_434_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_434_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_434_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_435_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_435_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_435_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_435_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_435_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_436_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_436_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_436_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_436_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_436_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_436_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_436_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_437_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_437_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_437_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_437_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_437_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_438_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_438_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_438_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_438_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_438_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_438_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_438_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_439_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_439_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_439_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_439_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_439_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_440_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_440_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_440_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_440_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_440_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_440_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_440_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_441_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_441_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_441_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_441_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_441_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_442_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_442_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_442_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_442_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_442_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_442_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_443_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_443_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_443_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_443_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_443_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_444_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_444_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_444_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_444_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_444_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_444_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_444_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_445_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_445_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_445_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_445_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_445_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_446_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_446_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_446_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_446_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_446_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_446_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_446_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_447_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_447_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_447_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_447_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_447_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_448_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_448_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_448_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_448_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_448_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_448_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_448_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_449_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_449_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_449_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_449_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_449_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_450_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_450_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_450_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_450_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_450_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_450_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_450_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_451_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_451_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_451_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_451_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_451_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_452_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_452_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_452_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_452_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_452_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_452_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_452_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_453_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_453_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_453_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_453_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_453_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_454_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_454_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_454_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_454_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_454_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_454_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_454_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_455_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_455_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_455_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_455_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_455_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_456_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_456_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_456_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_456_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_456_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_456_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_456_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_457_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_457_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_457_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_457_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_457_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_458_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_458_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_458_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_458_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_458_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_458_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_458_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_459_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_459_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_459_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_459_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_459_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_460_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_460_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_460_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_460_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_460_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_460_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_460_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_461_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_461_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_461_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_461_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_461_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_462_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_462_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_462_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_462_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_462_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_462_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_462_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_463_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_463_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_463_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_463_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_463_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_464_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_464_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_464_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_464_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_464_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_464_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_464_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_465_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_465_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_465_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_465_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_465_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_466_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_466_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_466_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_466_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_466_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_466_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_466_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_467_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_467_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_467_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_467_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_467_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_468_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_468_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_468_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_468_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_468_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_468_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_468_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_469_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_469_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_469_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_469_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_469_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_470_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_470_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_470_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_470_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_470_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_470_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_470_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_471_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_471_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_471_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_471_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_471_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_472_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_472_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_472_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_472_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_472_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_472_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_472_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_473_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_473_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_473_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_473_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_473_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_474_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_474_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_474_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_474_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_474_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_474_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_474_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_475_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_475_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_475_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_475_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_475_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_476_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_476_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_476_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_476_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_476_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_476_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_476_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_477_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_477_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_477_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_477_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_477_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_478_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_478_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_478_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_478_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_478_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_478_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_478_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_479_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_479_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_479_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_479_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_479_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_480_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_480_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_480_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_480_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_480_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_480_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_480_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_481_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_481_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_481_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_481_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_481_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_482_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_482_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_482_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_482_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_482_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_482_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_482_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_483_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_483_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_483_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_483_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_483_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_484_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_484_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_484_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_484_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_484_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_484_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_484_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_485_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_485_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_485_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_485_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_485_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_486_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_486_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_486_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_486_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_486_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_486_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_486_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_487_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_487_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_487_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_487_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_487_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_488_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_488_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_488_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_488_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_488_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_488_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_488_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_489_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_489_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_489_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_489_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_489_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_490_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_490_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_490_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_490_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_490_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_490_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_490_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_491_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_491_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_491_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_491_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_491_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_492_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_492_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_492_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_492_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_492_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_492_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_492_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_493_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_493_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_493_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_493_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_493_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_494_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_494_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_494_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_494_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_494_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_494_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_494_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_495_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_495_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_495_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_495_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_495_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_496_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_496_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_496_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_496_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_496_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_496_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_496_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_497_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_497_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_497_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_497_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_497_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_498_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_498_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_498_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_498_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_498_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_498_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_498_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_2458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_499_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_499_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_499_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_499_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_499_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_500_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_2636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_2668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_500_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_500_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_500_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_500_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_500_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_500_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_501_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_501_2370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_2374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_2454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_501_2486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_2490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_501_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_501_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_501_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_501_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_501_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_502_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_502_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_502_2364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_502_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_502_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_502_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_502_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_502_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_502_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_502_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_2330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_503_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_2366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_503_2368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_503_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_503_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_503_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_503_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_503_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_503_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_503_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_504_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_2280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_504_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_504_2336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_504_2346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_504_2373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_504_2383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_504_2410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_504_2416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_2635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_2667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_504_2669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_2928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_2992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_3024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_3348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_3380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_3704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_3736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_3996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_4060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_4092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_4416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_504_4448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_504_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_504_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_504_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_504_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_504_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_505_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_2314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_505_2342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_505_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_505_2362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_505_2479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_505_2487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_505_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_2814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_2846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_3170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_3202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_3526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_3558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_3882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_3914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_4238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_4270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_505_4466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_505_4530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_505_4562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_505_4566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_505_4568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_2298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_506_2348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_506_2356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_506_2358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_506_2411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_506_2477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_506_2485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_506_2489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_506_2491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_2654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_2832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_2914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_2978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_3156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_3334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_3512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_3690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_3868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_3900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_3982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_4046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_4078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_4096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_4160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_4224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_4256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_4274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_4338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_4402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_4434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_506_4452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_506_4516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_506_4548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_506_4564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_506_4568 ();
endmodule
