module parameterized_scrambler (clk,
    data_in,
    data_out,
    enable,
    rst_n,
    lfsr_state);
 input clk;
 input data_in;
 output data_out;
 input enable;
 input rst_n;
 output [7:0] lfsr_state;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire next_input;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _37_ (.A(rst_n),
    .Z(_08_));
 BUF_X2 _38_ (.A(enable),
    .Z(_09_));
 INV_X2 _39_ (.A(_09_),
    .ZN(_10_));
 NAND2_X1 _40_ (.A1(next_input),
    .A2(_10_),
    .ZN(_11_));
 NAND2_X1 _41_ (.A1(net4),
    .A2(_09_),
    .ZN(_12_));
 NAND3_X1 _42_ (.A1(_08_),
    .A2(_11_),
    .A3(_12_),
    .ZN(_00_));
 NAND2_X1 _43_ (.A1(net4),
    .A2(_10_),
    .ZN(_13_));
 NAND2_X1 _44_ (.A1(_09_),
    .A2(net5),
    .ZN(_14_));
 NAND3_X1 _45_ (.A1(_08_),
    .A2(_13_),
    .A3(_14_),
    .ZN(_01_));
 NAND2_X1 _46_ (.A1(_10_),
    .A2(net5),
    .ZN(_15_));
 NAND2_X1 _47_ (.A1(_09_),
    .A2(net6),
    .ZN(_16_));
 NAND3_X1 _48_ (.A1(_08_),
    .A2(_15_),
    .A3(_16_),
    .ZN(_02_));
 NAND2_X1 _49_ (.A1(net7),
    .A2(_09_),
    .ZN(_17_));
 NAND2_X1 _50_ (.A1(_10_),
    .A2(net6),
    .ZN(_18_));
 NAND3_X1 _51_ (.A1(_08_),
    .A2(_17_),
    .A3(_18_),
    .ZN(_03_));
 NAND2_X1 _52_ (.A1(net8),
    .A2(_09_),
    .ZN(_19_));
 NAND2_X1 _53_ (.A1(net7),
    .A2(_10_),
    .ZN(_20_));
 NAND3_X1 _54_ (.A1(_08_),
    .A2(_19_),
    .A3(_20_),
    .ZN(_04_));
 NAND2_X1 _55_ (.A1(net8),
    .A2(_10_),
    .ZN(_21_));
 NAND2_X1 _56_ (.A1(net9),
    .A2(_09_),
    .ZN(_22_));
 NAND3_X1 _57_ (.A1(_08_),
    .A2(_21_),
    .A3(_22_),
    .ZN(_05_));
 NAND2_X1 _58_ (.A1(net9),
    .A2(_10_),
    .ZN(_23_));
 NAND2_X1 _59_ (.A1(_09_),
    .A2(net10),
    .ZN(_24_));
 NAND3_X1 _60_ (.A1(_08_),
    .A2(_23_),
    .A3(_24_),
    .ZN(_06_));
 INV_X1 _61_ (.A(_08_),
    .ZN(_25_));
 AOI21_X1 _62_ (.A(_25_),
    .B1(net10),
    .B2(_10_),
    .ZN(_26_));
 XOR2_X1 _63_ (.A(net7),
    .B(net9),
    .Z(_27_));
 XNOR2_X1 _64_ (.A(net8),
    .B(_27_),
    .ZN(_28_));
 OAI21_X1 _65_ (.A(_26_),
    .B1(_28_),
    .B2(_10_),
    .ZN(_07_));
 XOR2_X1 _66_ (.A(next_input),
    .B(net1),
    .Z(net2));
 BUF_X1 _67_ (.A(next_input),
    .Z(net3));
 DFF_X1 \lfsr_reg[0]$_SDFFE_PN1P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(next_input),
    .QN(_36_));
 DFF_X1 \lfsr_reg[1]$_SDFFE_PN1P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_35_));
 DFF_X1 \lfsr_reg[2]$_SDFFE_PN1P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_34_));
 DFF_X1 \lfsr_reg[3]$_SDFFE_PN1P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net6),
    .QN(_33_));
 DFF_X2 \lfsr_reg[4]$_SDFFE_PN1P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net7),
    .QN(_32_));
 DFF_X2 \lfsr_reg[5]$_SDFFE_PN1P_  (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net8),
    .QN(_31_));
 DFF_X2 \lfsr_reg[6]$_SDFFE_PN1P_  (.D(_06_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net9),
    .QN(_30_));
 DFF_X1 \lfsr_reg[7]$_SDFFE_PN1P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_29_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_83 ();
 BUF_X1 input1 (.A(data_in),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(data_out));
 BUF_X1 output3 (.A(net3),
    .Z(lfsr_state[0]));
 BUF_X1 output4 (.A(net4),
    .Z(lfsr_state[1]));
 BUF_X1 output5 (.A(net5),
    .Z(lfsr_state[2]));
 BUF_X1 output6 (.A(net6),
    .Z(lfsr_state[3]));
 BUF_X1 output7 (.A(net7),
    .Z(lfsr_state[4]));
 BUF_X1 output8 (.A(net8),
    .Z(lfsr_state[5]));
 BUF_X1 output9 (.A(net9),
    .Z(lfsr_state[6]));
 BUF_X1 output10 (.A(net10),
    .Z(lfsr_state[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_129 ();
 FILLCELL_X2 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_147 ();
 FILLCELL_X4 FILLER_0_151 ();
 FILLCELL_X2 FILLER_0_155 ();
 FILLCELL_X32 FILLER_0_160 ();
 FILLCELL_X32 FILLER_0_192 ();
 FILLCELL_X32 FILLER_0_224 ();
 FILLCELL_X32 FILLER_0_256 ();
 FILLCELL_X16 FILLER_0_288 ();
 FILLCELL_X8 FILLER_0_304 ();
 FILLCELL_X2 FILLER_0_312 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_145 ();
 FILLCELL_X2 FILLER_1_149 ();
 FILLCELL_X1 FILLER_1_151 ();
 FILLCELL_X32 FILLER_1_155 ();
 FILLCELL_X32 FILLER_1_187 ();
 FILLCELL_X32 FILLER_1_219 ();
 FILLCELL_X32 FILLER_1_251 ();
 FILLCELL_X16 FILLER_1_283 ();
 FILLCELL_X8 FILLER_1_299 ();
 FILLCELL_X4 FILLER_1_307 ();
 FILLCELL_X2 FILLER_1_311 ();
 FILLCELL_X1 FILLER_1_313 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X16 FILLER_2_289 ();
 FILLCELL_X8 FILLER_2_305 ();
 FILLCELL_X1 FILLER_2_313 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X16 FILLER_3_289 ();
 FILLCELL_X8 FILLER_3_305 ();
 FILLCELL_X1 FILLER_3_313 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X16 FILLER_4_289 ();
 FILLCELL_X8 FILLER_4_305 ();
 FILLCELL_X1 FILLER_4_313 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X16 FILLER_5_289 ();
 FILLCELL_X8 FILLER_5_305 ();
 FILLCELL_X1 FILLER_5_313 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X16 FILLER_6_289 ();
 FILLCELL_X8 FILLER_6_305 ();
 FILLCELL_X1 FILLER_6_313 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X16 FILLER_7_289 ();
 FILLCELL_X8 FILLER_7_305 ();
 FILLCELL_X1 FILLER_7_313 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X16 FILLER_8_289 ();
 FILLCELL_X8 FILLER_8_305 ();
 FILLCELL_X1 FILLER_8_313 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X16 FILLER_9_289 ();
 FILLCELL_X8 FILLER_9_305 ();
 FILLCELL_X1 FILLER_9_313 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X16 FILLER_10_289 ();
 FILLCELL_X8 FILLER_10_305 ();
 FILLCELL_X1 FILLER_10_313 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X16 FILLER_11_289 ();
 FILLCELL_X8 FILLER_11_305 ();
 FILLCELL_X1 FILLER_11_313 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X16 FILLER_12_289 ();
 FILLCELL_X8 FILLER_12_305 ();
 FILLCELL_X1 FILLER_12_313 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X16 FILLER_13_289 ();
 FILLCELL_X8 FILLER_13_305 ();
 FILLCELL_X1 FILLER_13_313 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X16 FILLER_14_289 ();
 FILLCELL_X8 FILLER_14_305 ();
 FILLCELL_X1 FILLER_14_313 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X16 FILLER_15_289 ();
 FILLCELL_X8 FILLER_15_305 ();
 FILLCELL_X1 FILLER_15_313 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X16 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_145 ();
 FILLCELL_X1 FILLER_16_153 ();
 FILLCELL_X8 FILLER_16_160 ();
 FILLCELL_X32 FILLER_16_171 ();
 FILLCELL_X32 FILLER_16_203 ();
 FILLCELL_X32 FILLER_16_235 ();
 FILLCELL_X32 FILLER_16_267 ();
 FILLCELL_X8 FILLER_16_299 ();
 FILLCELL_X4 FILLER_16_307 ();
 FILLCELL_X2 FILLER_16_311 ();
 FILLCELL_X1 FILLER_16_313 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_137 ();
 FILLCELL_X1 FILLER_17_141 ();
 FILLCELL_X1 FILLER_17_165 ();
 FILLCELL_X32 FILLER_17_190 ();
 FILLCELL_X32 FILLER_17_222 ();
 FILLCELL_X16 FILLER_17_254 ();
 FILLCELL_X4 FILLER_17_270 ();
 FILLCELL_X2 FILLER_17_274 ();
 FILLCELL_X32 FILLER_17_279 ();
 FILLCELL_X2 FILLER_17_311 ();
 FILLCELL_X1 FILLER_17_313 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X16 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_145 ();
 FILLCELL_X1 FILLER_18_163 ();
 FILLCELL_X1 FILLER_18_167 ();
 FILLCELL_X4 FILLER_18_172 ();
 FILLCELL_X32 FILLER_18_208 ();
 FILLCELL_X32 FILLER_18_240 ();
 FILLCELL_X32 FILLER_18_272 ();
 FILLCELL_X8 FILLER_18_304 ();
 FILLCELL_X2 FILLER_18_312 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X16 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_145 ();
 FILLCELL_X4 FILLER_19_153 ();
 FILLCELL_X1 FILLER_19_157 ();
 FILLCELL_X32 FILLER_19_164 ();
 FILLCELL_X32 FILLER_19_196 ();
 FILLCELL_X32 FILLER_19_228 ();
 FILLCELL_X32 FILLER_19_260 ();
 FILLCELL_X16 FILLER_19_292 ();
 FILLCELL_X4 FILLER_19_308 ();
 FILLCELL_X2 FILLER_19_312 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X8 FILLER_20_129 ();
 FILLCELL_X4 FILLER_20_137 ();
 FILLCELL_X1 FILLER_20_141 ();
 FILLCELL_X16 FILLER_20_165 ();
 FILLCELL_X8 FILLER_20_181 ();
 FILLCELL_X2 FILLER_20_189 ();
 FILLCELL_X1 FILLER_20_191 ();
 FILLCELL_X32 FILLER_20_196 ();
 FILLCELL_X32 FILLER_20_228 ();
 FILLCELL_X32 FILLER_20_260 ();
 FILLCELL_X16 FILLER_20_292 ();
 FILLCELL_X4 FILLER_20_308 ();
 FILLCELL_X2 FILLER_20_312 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X16 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_145 ();
 FILLCELL_X16 FILLER_21_156 ();
 FILLCELL_X4 FILLER_21_172 ();
 FILLCELL_X2 FILLER_21_176 ();
 FILLCELL_X1 FILLER_21_178 ();
 FILLCELL_X32 FILLER_21_182 ();
 FILLCELL_X32 FILLER_21_214 ();
 FILLCELL_X32 FILLER_21_246 ();
 FILLCELL_X32 FILLER_21_278 ();
 FILLCELL_X4 FILLER_21_310 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X16 FILLER_22_129 ();
 FILLCELL_X4 FILLER_22_145 ();
 FILLCELL_X2 FILLER_22_149 ();
 FILLCELL_X16 FILLER_22_158 ();
 FILLCELL_X32 FILLER_22_179 ();
 FILLCELL_X32 FILLER_22_211 ();
 FILLCELL_X32 FILLER_22_243 ();
 FILLCELL_X32 FILLER_22_275 ();
 FILLCELL_X4 FILLER_22_307 ();
 FILLCELL_X2 FILLER_22_311 ();
 FILLCELL_X1 FILLER_22_313 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X8 FILLER_23_129 ();
 FILLCELL_X2 FILLER_23_137 ();
 FILLCELL_X1 FILLER_23_139 ();
 FILLCELL_X16 FILLER_23_157 ();
 FILLCELL_X2 FILLER_23_173 ();
 FILLCELL_X1 FILLER_23_175 ();
 FILLCELL_X2 FILLER_23_183 ();
 FILLCELL_X32 FILLER_23_195 ();
 FILLCELL_X32 FILLER_23_227 ();
 FILLCELL_X32 FILLER_23_259 ();
 FILLCELL_X8 FILLER_23_291 ();
 FILLCELL_X4 FILLER_23_299 ();
 FILLCELL_X2 FILLER_23_303 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X4 FILLER_24_145 ();
 FILLCELL_X1 FILLER_24_149 ();
 FILLCELL_X8 FILLER_24_160 ();
 FILLCELL_X2 FILLER_24_168 ();
 FILLCELL_X1 FILLER_24_170 ();
 FILLCELL_X32 FILLER_24_208 ();
 FILLCELL_X32 FILLER_24_240 ();
 FILLCELL_X16 FILLER_24_272 ();
 FILLCELL_X8 FILLER_24_288 ();
 FILLCELL_X4 FILLER_24_296 ();
 FILLCELL_X2 FILLER_24_300 ();
 FILLCELL_X2 FILLER_24_305 ();
 FILLCELL_X1 FILLER_24_307 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X16 FILLER_25_129 ();
 FILLCELL_X4 FILLER_25_145 ();
 FILLCELL_X2 FILLER_25_149 ();
 FILLCELL_X1 FILLER_25_151 ();
 FILLCELL_X32 FILLER_25_169 ();
 FILLCELL_X32 FILLER_25_201 ();
 FILLCELL_X32 FILLER_25_233 ();
 FILLCELL_X32 FILLER_25_265 ();
 FILLCELL_X16 FILLER_25_297 ();
 FILLCELL_X1 FILLER_25_313 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X4 FILLER_26_161 ();
 FILLCELL_X2 FILLER_26_165 ();
 FILLCELL_X1 FILLER_26_167 ();
 FILLCELL_X32 FILLER_26_177 ();
 FILLCELL_X32 FILLER_26_209 ();
 FILLCELL_X32 FILLER_26_241 ();
 FILLCELL_X32 FILLER_26_273 ();
 FILLCELL_X8 FILLER_26_305 ();
 FILLCELL_X1 FILLER_26_313 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X16 FILLER_27_289 ();
 FILLCELL_X8 FILLER_27_305 ();
 FILLCELL_X1 FILLER_27_313 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X16 FILLER_28_289 ();
 FILLCELL_X8 FILLER_28_305 ();
 FILLCELL_X1 FILLER_28_313 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X16 FILLER_29_289 ();
 FILLCELL_X8 FILLER_29_305 ();
 FILLCELL_X1 FILLER_29_313 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X16 FILLER_30_289 ();
 FILLCELL_X8 FILLER_30_305 ();
 FILLCELL_X1 FILLER_30_313 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X16 FILLER_31_289 ();
 FILLCELL_X8 FILLER_31_305 ();
 FILLCELL_X1 FILLER_31_313 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X16 FILLER_32_289 ();
 FILLCELL_X8 FILLER_32_305 ();
 FILLCELL_X1 FILLER_32_313 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X16 FILLER_33_289 ();
 FILLCELL_X8 FILLER_33_305 ();
 FILLCELL_X1 FILLER_33_313 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X16 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_305 ();
 FILLCELL_X1 FILLER_34_313 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X16 FILLER_35_289 ();
 FILLCELL_X8 FILLER_35_305 ();
 FILLCELL_X1 FILLER_35_313 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X16 FILLER_36_289 ();
 FILLCELL_X8 FILLER_36_305 ();
 FILLCELL_X1 FILLER_36_313 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X16 FILLER_37_289 ();
 FILLCELL_X8 FILLER_37_305 ();
 FILLCELL_X1 FILLER_37_313 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X16 FILLER_38_289 ();
 FILLCELL_X8 FILLER_38_305 ();
 FILLCELL_X1 FILLER_38_313 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X16 FILLER_39_289 ();
 FILLCELL_X8 FILLER_39_305 ();
 FILLCELL_X1 FILLER_39_313 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X16 FILLER_40_289 ();
 FILLCELL_X8 FILLER_40_305 ();
 FILLCELL_X1 FILLER_40_313 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X16 FILLER_41_129 ();
 FILLCELL_X8 FILLER_41_148 ();
 FILLCELL_X1 FILLER_41_156 ();
 FILLCELL_X16 FILLER_41_160 ();
 FILLCELL_X4 FILLER_41_176 ();
 FILLCELL_X1 FILLER_41_180 ();
 FILLCELL_X32 FILLER_41_184 ();
 FILLCELL_X32 FILLER_41_216 ();
 FILLCELL_X32 FILLER_41_248 ();
 FILLCELL_X32 FILLER_41_280 ();
 FILLCELL_X2 FILLER_41_312 ();
endmodule
