module cordic_core (x_in,
    x_out,
    y_in,
    y_out,
    z_in);
 input [15:0] x_in;
 output [15:0] x_out;
 input [15:0] y_in;
 output [15:0] y_out;
 input [15:0] z_in;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire net2;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire net1;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net197;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net228;
 wire net229;
 wire net233;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net173;
 wire net174;
 wire net175;
 wire net180;
 wire net181;
 wire net195;
 wire net196;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net264;
 wire net272;

 sky130_fd_sc_hd__inv_1 _3747_ (.A(net68),
    .Y(_3684_));
 sky130_fd_sc_hd__nor3_1 _3748_ (.A(net70),
    .B(net69),
    .C(net62),
    .Y(_0000_));
 sky130_fd_sc_hd__nor4_2 _3749_ (.A(net74),
    .B(net73),
    .C(net72),
    .D(net71),
    .Y(_0001_));
 sky130_fd_sc_hd__and2_0 _3750_ (.A(_0000_),
    .B(_0001_),
    .X(_0002_));
 sky130_fd_sc_hd__nor4_2 _3751_ (.A(net66),
    .B(net65),
    .C(net64),
    .D(net63),
    .Y(_0003_));
 sky130_fd_sc_hd__and2b_2 _3752_ (.A_N(_3687_),
    .B(net68),
    .X(_0004_));
 sky130_fd_sc_hd__or3_4 _3753_ (.A(net77),
    .B(net76),
    .C(net75),
    .X(_0005_));
 sky130_fd_sc_hd__nor4_4 _3754_ (.A(_0004_),
    .B(_3685_),
    .C(net67),
    .D(_0005_),
    .Y(_0006_));
 sky130_fd_sc_hd__a32o_4 _3755_ (.A1(_0006_),
    .A2(_0003_),
    .A3(_0002_),
    .B1(_3685_),
    .B2(net68),
    .X(_0007_));
 sky130_fd_sc_hd__inv_6 _3756_ (.A(_0007_),
    .Y(_0008_));
 sky130_fd_sc_hd__buf_8 _3757_ (.A(_0008_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_12 _3758_ (.A(_0009_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_8 _3759_ (.A(_0010_),
    .X(_2091_));
 sky130_fd_sc_hd__nand2_1 _3760_ (.A(_2081_),
    .B(_2091_),
    .Y(_0011_));
 sky130_fd_sc_hd__buf_4 _3761_ (.A(_0007_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_4 _3762_ (.A(_0012_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _3763_ (.A(_0013_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _3764_ (.A(_0014_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _3765_ (.A(_0015_),
    .X(_0016_));
 sky130_fd_sc_hd__nand2_1 _3766_ (.A(_2085_),
    .B(_0016_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _3767_ (.A(_0011_),
    .B(_0017_),
    .Y(_2207_));
 sky130_fd_sc_hd__inv_1 _3768_ (.A(_2207_),
    .Y(_2096_));
 sky130_fd_sc_hd__nor2b_1 _3769_ (.A(_2086_),
    .B_N(_2201_),
    .Y(_0018_));
 sky130_fd_sc_hd__clkbuf_2 _3770_ (.A(_2219_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _3771_ (.A(_2211_),
    .X(_0020_));
 sky130_fd_sc_hd__o21a_1 _3772_ (.A1(_0019_),
    .A2(_2218_),
    .B1(_0020_),
    .X(_0021_));
 sky130_fd_sc_hd__o31a_2 _3773_ (.A1(_2202_),
    .A2(_2218_),
    .A3(_0018_),
    .B1(_0021_),
    .X(_0022_));
 sky130_fd_sc_hd__o21a_1 _3774_ (.A1(_2202_),
    .A2(_0018_),
    .B1(_0019_),
    .X(_0023_));
 sky130_fd_sc_hd__nor3_1 _3775_ (.A(_0020_),
    .B(_2218_),
    .C(_0023_),
    .Y(_0024_));
 sky130_fd_sc_hd__nor2_1 _3776_ (.A(_0022_),
    .B(_0024_),
    .Y(_0025_));
 sky130_fd_sc_hd__nor3b_1 _3777_ (.A(_0019_),
    .B(_2201_),
    .C_N(_2199_),
    .Y(_0026_));
 sky130_fd_sc_hd__nor2b_1 _3778_ (.A(_0019_),
    .B_N(_2205_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor3_1 _3779_ (.A(_2223_),
    .B(_0026_),
    .C(_0027_),
    .Y(_0028_));
 sky130_fd_sc_hd__xnor2_2 _3780_ (.A(_0020_),
    .B(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_1 _3781_ (.A(_0015_),
    .B(_0029_),
    .Y(_0030_));
 sky130_fd_sc_hd__a21oi_1 _3782_ (.A1(_0015_),
    .A2(_0025_),
    .B1(_0030_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_1 _3783_ (.A(_0031_),
    .Y(_2272_));
 sky130_fd_sc_hd__clkbuf_4 _3784_ (.A(_0019_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_2 _3785_ (.A(_2084_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _3786_ (.A(_2087_),
    .B(_0014_),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_0 _3787_ (.A1(_0033_),
    .A2(_0014_),
    .B1(_0034_),
    .Y(_0035_));
 sky130_fd_sc_hd__xnor2_1 _3788_ (.A(_0032_),
    .B(_0035_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_1 _3789_ (.A(_2085_),
    .B(_2091_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _3790_ (.A(_2088_),
    .B(_0016_),
    .Y(_0037_));
 sky130_fd_sc_hd__nand2_2 _3791_ (.A(_0036_),
    .B(_0037_),
    .Y(_2101_));
 sky130_fd_sc_hd__inv_1 _3792_ (.A(_2101_),
    .Y(_2105_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(net67),
    .Y(_3683_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(_0000_),
    .B(_0001_),
    .Y(_0038_));
 sky130_fd_sc_hd__or2_0 _3795_ (.A(_0038_),
    .B(_0005_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_1 _3796_ (.A(_3685_),
    .B(_0004_),
    .Y(_0040_));
 sky130_fd_sc_hd__buf_2 _3797_ (.A(_0040_),
    .X(_0041_));
 sky130_fd_sc_hd__o41ai_2 _3798_ (.A1(net65),
    .A2(net64),
    .A3(net63),
    .A4(_0039_),
    .B1(_0041_),
    .Y(_0042_));
 sky130_fd_sc_hd__xnor2_2 _3799_ (.A(net66),
    .B(_0042_),
    .Y(_2089_));
 sky130_fd_sc_hd__inv_1 _3800_ (.A(_2089_),
    .Y(_2284_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_0033_),
    .B(_0015_),
    .Y(_0043_));
 sky130_fd_sc_hd__o21ai_1 _3802_ (.A1(_2080_),
    .A2(_0015_),
    .B1(_0043_),
    .Y(_0044_));
 sky130_fd_sc_hd__xnor2_2 _3803_ (.A(_0032_),
    .B(_0044_),
    .Y(_2279_));
 sky130_fd_sc_hd__inv_1 _3804_ (.A(_2279_),
    .Y(_2227_));
 sky130_fd_sc_hd__inv_1 _3805_ (.A(_2276_),
    .Y(_2231_));
 sky130_fd_sc_hd__buf_12 _3806_ (.A(_2092_),
    .X(_0045_));
 sky130_fd_sc_hd__clkinv_8 _3807_ (.A(_0045_),
    .Y(_2111_));
 sky130_fd_sc_hd__mux2_1 _3808_ (.A0(_2233_),
    .A1(_2276_),
    .S(_2111_),
    .X(_2234_));
 sky130_fd_sc_hd__inv_1 _3809_ (.A(_2234_),
    .Y(_2095_));
 sky130_fd_sc_hd__xnor2_2 _3810_ (.A(_2230_),
    .B(_2097_),
    .Y(_2237_));
 sky130_fd_sc_hd__inv_1 _3811_ (.A(_2237_),
    .Y(_2428_));
 sky130_fd_sc_hd__clkbuf_4 _3812_ (.A(_2241_),
    .X(_0046_));
 sky130_fd_sc_hd__clkinvlp_4 _3813_ (.A(_0046_),
    .Y(_0047_));
 sky130_fd_sc_hd__nor2b_1 _3814_ (.A(_0046_),
    .B_N(_2249_),
    .Y(_0048_));
 sky130_fd_sc_hd__o21a_1 _3815_ (.A1(_2210_),
    .A2(_0022_),
    .B1(_0048_),
    .X(_0049_));
 sky130_fd_sc_hd__nor4_1 _3816_ (.A(_0047_),
    .B(_2210_),
    .C(_2248_),
    .D(_0022_),
    .Y(_0050_));
 sky130_fd_sc_hd__buf_4 _3817_ (.A(_2249_),
    .X(_0051_));
 sky130_fd_sc_hd__nor3_1 _3818_ (.A(_0051_),
    .B(_0047_),
    .C(_2248_),
    .Y(_0052_));
 sky130_fd_sc_hd__a2111oi_4 _3819_ (.A1(_0047_),
    .A2(_2248_),
    .B1(_0049_),
    .C1(_0050_),
    .D1(_0052_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_1 _3820_ (.A(_0020_),
    .Y(_0054_));
 sky130_fd_sc_hd__o31a_2 _3821_ (.A1(_2223_),
    .A2(_0026_),
    .A3(_0027_),
    .B1(_0054_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2b_1 _3822_ (.A_N(_2215_),
    .B(_0046_),
    .Y(_0056_));
 sky130_fd_sc_hd__buf_2 _3823_ (.A(_0046_),
    .X(_0057_));
 sky130_fd_sc_hd__nor2_1 _3824_ (.A(_0051_),
    .B(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__o311ai_1 _3825_ (.A1(_2223_),
    .A2(_0026_),
    .A3(_0027_),
    .B1(_0058_),
    .C1(_0054_),
    .Y(_0059_));
 sky130_fd_sc_hd__nor2b_1 _3826_ (.A(_2249_),
    .B_N(_2215_),
    .Y(_0060_));
 sky130_fd_sc_hd__and3b_1 _3827_ (.A_N(_2253_),
    .B(_0057_),
    .C(_0051_),
    .X(_0061_));
 sky130_fd_sc_hd__nor2b_1 _3828_ (.A(_0046_),
    .B_N(_2253_),
    .Y(_0062_));
 sky130_fd_sc_hd__a211oi_1 _3829_ (.A1(_0047_),
    .A2(_0060_),
    .B1(_0061_),
    .C1(_0062_),
    .Y(_0063_));
 sky130_fd_sc_hd__o311a_2 _3830_ (.A1(_2253_),
    .A2(_0055_),
    .A3(_0056_),
    .B1(_0059_),
    .C1(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(net172),
    .B(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__o21ai_2 _3832_ (.A1(net172),
    .A2(_0053_),
    .B1(_0065_),
    .Y(_2264_));
 sky130_fd_sc_hd__buf_2 _3833_ (.A(_2257_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_0 _3834_ (.A(_2251_),
    .B(_2243_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2b_1 _3835_ (.A(_2080_),
    .B_N(_0019_),
    .Y(_0068_));
 sky130_fd_sc_hd__o21a_1 _3836_ (.A1(_0020_),
    .A2(_2213_),
    .B1(_0051_),
    .X(_0069_));
 sky130_fd_sc_hd__o31a_2 _3837_ (.A1(_2221_),
    .A2(_2213_),
    .A3(_0068_),
    .B1(_0069_),
    .X(_0070_));
 sky130_fd_sc_hd__o22a_1 _3838_ (.A1(_0057_),
    .A2(_2243_),
    .B1(_0067_),
    .B2(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__xnor2_1 _3839_ (.A(_0066_),
    .B(_0071_),
    .Y(_0072_));
 sky130_fd_sc_hd__clkinvlp_4 _3840_ (.A(_2257_),
    .Y(_0073_));
 sky130_fd_sc_hd__o21bai_1 _3841_ (.A1(_0019_),
    .A2(_0033_),
    .B1_N(_2223_),
    .Y(_0074_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(_0020_),
    .B(_2249_),
    .Y(_0075_));
 sky130_fd_sc_hd__a211o_1 _3843_ (.A1(_0074_),
    .A2(_0075_),
    .B1(_2253_),
    .C1(_0060_),
    .X(_0076_));
 sky130_fd_sc_hd__a21oi_1 _3844_ (.A1(_0047_),
    .A2(_0076_),
    .B1(_2245_),
    .Y(_0077_));
 sky130_fd_sc_hd__xnor2_2 _3845_ (.A(_0073_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor2_1 _3846_ (.A(_0010_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__a21oi_2 _3847_ (.A1(_0010_),
    .A2(_0072_),
    .B1(_0079_),
    .Y(_2392_));
 sky130_fd_sc_hd__nor2b_2 _3848_ (.A(_2079_),
    .B_N(_2201_),
    .Y(_0080_));
 sky130_fd_sc_hd__o21a_1 _3849_ (.A1(_0019_),
    .A2(_2221_),
    .B1(_0020_),
    .X(_0081_));
 sky130_fd_sc_hd__o31a_1 _3850_ (.A1(_2221_),
    .A2(_2203_),
    .A3(_0080_),
    .B1(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2b_1 _3851_ (.A_N(_2251_),
    .B(_0057_),
    .Y(_0083_));
 sky130_fd_sc_hd__o311ai_1 _3852_ (.A1(_2221_),
    .A2(_2203_),
    .A3(_0080_),
    .B1(_0081_),
    .C1(_0048_),
    .Y(_0084_));
 sky130_fd_sc_hd__nor3b_1 _3853_ (.A(_0051_),
    .B(_2251_),
    .C_N(_0057_),
    .Y(_0085_));
 sky130_fd_sc_hd__a221oi_1 _3854_ (.A1(_0047_),
    .A2(_2251_),
    .B1(_2213_),
    .B2(_0048_),
    .C1(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__o311ai_2 _3855_ (.A1(_2213_),
    .A2(_0082_),
    .A3(_0083_),
    .B1(_0084_),
    .C1(_0086_),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2b_1 _3856_ (.A_N(_0064_),
    .B(_0013_),
    .Y(_0088_));
 sky130_fd_sc_hd__o21a_1 _3857_ (.A1(_0014_),
    .A2(_0087_),
    .B1(_0088_),
    .X(_2396_));
 sky130_fd_sc_hd__a21oi_1 _3858_ (.A1(_0054_),
    .A2(_0074_),
    .B1(_2215_),
    .Y(_0089_));
 sky130_fd_sc_hd__xnor2_2 _3859_ (.A(_0051_),
    .B(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_0 _3860_ (.A1(_2221_),
    .A2(_0068_),
    .B1(_0020_),
    .Y(_0091_));
 sky130_fd_sc_hd__nor2_1 _3861_ (.A(_0051_),
    .B(_2213_),
    .Y(_0092_));
 sky130_fd_sc_hd__a21oi_1 _3862_ (.A1(_0091_),
    .A2(_0092_),
    .B1(_0070_),
    .Y(_0093_));
 sky130_fd_sc_hd__nor2_1 _3863_ (.A(_0016_),
    .B(_0093_),
    .Y(_0094_));
 sky130_fd_sc_hd__a21oi_2 _3864_ (.A1(_0016_),
    .A2(_0090_),
    .B1(_0094_),
    .Y(_2400_));
 sky130_fd_sc_hd__o31ai_4 _3865_ (.A1(_2221_),
    .A2(_2203_),
    .A3(_0080_),
    .B1(_0081_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_1 _3866_ (.A(_2221_),
    .Y(_0096_));
 sky130_fd_sc_hd__o21ai_0 _3867_ (.A1(_2203_),
    .A2(_0080_),
    .B1(_0032_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand3_1 _3868_ (.A(_0054_),
    .B(_0096_),
    .C(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__a21oi_1 _3869_ (.A1(_0095_),
    .A2(_0098_),
    .B1(_0014_),
    .Y(_0099_));
 sky130_fd_sc_hd__a21oi_2 _3870_ (.A1(_0015_),
    .A2(_0029_),
    .B1(_0099_),
    .Y(_2317_));
 sky130_fd_sc_hd__xnor2_1 _3871_ (.A(_0032_),
    .B(_2080_),
    .Y(_0100_));
 sky130_fd_sc_hd__nor2_1 _3872_ (.A(_2081_),
    .B(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__a2111oi_0 _3873_ (.A1(_0095_),
    .A2(_0098_),
    .B1(_0087_),
    .C1(_0013_),
    .D1(_0093_),
    .Y(_0102_));
 sky130_fd_sc_hd__xor2_1 _3874_ (.A(_0032_),
    .B(_0033_),
    .X(_0103_));
 sky130_fd_sc_hd__nor2_1 _3875_ (.A(_2085_),
    .B(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand3_1 _3876_ (.A(_0029_),
    .B(_0090_),
    .C(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__o2bb2ai_1 _3877_ (.A1_N(_0101_),
    .A2_N(_0102_),
    .B1(_0105_),
    .B2(_0088_),
    .Y(_0106_));
 sky130_fd_sc_hd__nor2_1 _3878_ (.A(net16),
    .B(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__xnor2_1 _3879_ (.A(_2392_),
    .B(_0107_),
    .Y(_2263_));
 sky130_fd_sc_hd__nor2b_1 _3880_ (.A(_2087_),
    .B_N(_0019_),
    .Y(_0108_));
 sky130_fd_sc_hd__o21ai_0 _3881_ (.A1(_2218_),
    .A2(_0108_),
    .B1(_0020_),
    .Y(_0109_));
 sky130_fd_sc_hd__nor2_1 _3882_ (.A(_0051_),
    .B(_2210_),
    .Y(_0110_));
 sky130_fd_sc_hd__o21a_1 _3883_ (.A1(_0020_),
    .A2(_2210_),
    .B1(_2249_),
    .X(_0111_));
 sky130_fd_sc_hd__o31a_2 _3884_ (.A1(_2218_),
    .A2(_2210_),
    .A3(_0108_),
    .B1(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__a21oi_1 _3885_ (.A1(_0109_),
    .A2(_0110_),
    .B1(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__nand2_1 _3886_ (.A(_0016_),
    .B(_0113_),
    .Y(_0114_));
 sky130_fd_sc_hd__o21ai_1 _3887_ (.A1(_0015_),
    .A2(_0090_),
    .B1(_0114_),
    .Y(_2268_));
 sky130_fd_sc_hd__buf_2 _3888_ (.A(_0045_),
    .X(_0115_));
 sky130_fd_sc_hd__a211oi_1 _3889_ (.A1(_0095_),
    .A2(_0098_),
    .B1(_0093_),
    .C1(_0014_),
    .Y(_0116_));
 sky130_fd_sc_hd__and3_1 _3890_ (.A(_0013_),
    .B(_0029_),
    .C(_0090_),
    .X(_0117_));
 sky130_fd_sc_hd__o21ai_1 _3891_ (.A1(_0116_),
    .A2(_0117_),
    .B1(_2280_),
    .Y(_0118_));
 sky130_fd_sc_hd__nand2_1 _3892_ (.A(_0115_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__xor2_1 _3893_ (.A(_2396_),
    .B(_0119_),
    .X(_2267_));
 sky130_fd_sc_hd__nand3b_1 _3894_ (.A_N(_2085_),
    .B(_0033_),
    .C(_0014_),
    .Y(_0120_));
 sky130_fd_sc_hd__o311a_1 _3895_ (.A1(_2081_),
    .A2(_2080_),
    .A3(_0014_),
    .B1(_0120_),
    .C1(_0032_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _3896_ (.A(_2081_),
    .B(_0015_),
    .Y(_0122_));
 sky130_fd_sc_hd__nor3_1 _3897_ (.A(_2085_),
    .B(_0033_),
    .C(net172),
    .Y(_0123_));
 sky130_fd_sc_hd__a211oi_1 _3898_ (.A1(_2080_),
    .A2(_0122_),
    .B1(_0123_),
    .C1(_0032_),
    .Y(_0124_));
 sky130_fd_sc_hd__buf_2 _3899_ (.A(_0045_),
    .X(_0125_));
 sky130_fd_sc_hd__o31ai_1 _3900_ (.A1(_2317_),
    .A2(_0121_),
    .A3(_0124_),
    .B1(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__xor2_1 _3901_ (.A(_2400_),
    .B(_0126_),
    .X(_2271_));
 sky130_fd_sc_hd__nor2_1 _3902_ (.A(_2111_),
    .B(_2280_),
    .Y(_0127_));
 sky130_fd_sc_hd__xnor2_1 _3903_ (.A(_2317_),
    .B(_0127_),
    .Y(_2275_));
 sky130_fd_sc_hd__nor2_1 _3904_ (.A(_0115_),
    .B(_2279_),
    .Y(_0128_));
 sky130_fd_sc_hd__a21oi_2 _3905_ (.A1(_0115_),
    .A2(_2281_),
    .B1(_0128_),
    .Y(_2100_));
 sky130_fd_sc_hd__inv_1 _3906_ (.A(_2104_),
    .Y(_2099_));
 sky130_fd_sc_hd__nor2b_1 _3907_ (.A(_2104_),
    .B_N(_2283_),
    .Y(_0129_));
 sky130_fd_sc_hd__o21ai_0 _3908_ (.A1(_2282_),
    .A2(_0129_),
    .B1(_2278_),
    .Y(_0130_));
 sky130_fd_sc_hd__nor2_1 _3909_ (.A(_2274_),
    .B(_2277_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21a_1 _3910_ (.A1(_2278_),
    .A2(_2277_),
    .B1(_2274_),
    .X(_0132_));
 sky130_fd_sc_hd__o31a_1 _3911_ (.A1(_2277_),
    .A2(_2282_),
    .A3(_0129_),
    .B1(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a21oi_2 _3912_ (.A1(_0130_),
    .A2(_0131_),
    .B1(_0133_),
    .Y(_2420_));
 sky130_fd_sc_hd__inv_1 _3913_ (.A(_2420_),
    .Y(_2328_));
 sky130_fd_sc_hd__xor2_2 _3914_ (.A(_2278_),
    .B(_2102_),
    .X(_2424_));
 sky130_fd_sc_hd__inv_1 _3915_ (.A(_2424_),
    .Y(_2327_));
 sky130_fd_sc_hd__o21ai_0 _3916_ (.A1(_2273_),
    .A2(_0133_),
    .B1(_2270_),
    .Y(_0134_));
 sky130_fd_sc_hd__nor2_1 _3917_ (.A(_2266_),
    .B(_2269_),
    .Y(_0135_));
 sky130_fd_sc_hd__o21a_1 _3918_ (.A1(_2270_),
    .A2(_2269_),
    .B1(_2266_),
    .X(_0136_));
 sky130_fd_sc_hd__o31a_1 _3919_ (.A1(_2269_),
    .A2(_2273_),
    .A3(_0133_),
    .B1(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__a21oi_2 _3920_ (.A1(_0134_),
    .A2(_0135_),
    .B1(_0137_),
    .Y(_2412_));
 sky130_fd_sc_hd__buf_8 _3921_ (.A(net62),
    .X(_0138_));
 sky130_fd_sc_hd__clkinv_8 _3922_ (.A(_0138_),
    .Y(_2122_));
 sky130_fd_sc_hd__o31a_1 _3923_ (.A1(_2472_),
    .A2(_3685_),
    .A3(_0004_),
    .B1(net70),
    .X(_0139_));
 sky130_fd_sc_hd__nor4_1 _3924_ (.A(net70),
    .B(_2472_),
    .C(_3685_),
    .D(_0004_),
    .Y(_0140_));
 sky130_fd_sc_hd__nor2_1 _3925_ (.A(_0139_),
    .B(_0140_),
    .Y(_2110_));
 sky130_fd_sc_hd__inv_1 _3926_ (.A(_2294_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21oi_2 _3927_ (.A1(_2313_),
    .A2(_2314_),
    .B1(_2312_),
    .Y(_0142_));
 sky130_fd_sc_hd__o211ai_1 _3928_ (.A1(_0139_),
    .A2(_0140_),
    .B1(_2313_),
    .C1(_2315_),
    .Y(_0143_));
 sky130_fd_sc_hd__a21boi_4 _3929_ (.A1(_0143_),
    .A2(_0142_),
    .B1_N(_2310_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_1 _3930_ (.A(_2307_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_1 _3931_ (.A(_2301_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand2_1 _3932_ (.A(_2298_),
    .B(_2304_),
    .Y(_0147_));
 sky130_fd_sc_hd__nor3_2 _3933_ (.A(_0145_),
    .B(_0146_),
    .C(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__o21ai_4 _3934_ (.A1(_0144_),
    .A2(_2309_),
    .B1(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__a21oi_2 _3935_ (.A1(_2304_),
    .A2(_2306_),
    .B1(_2303_),
    .Y(_0150_));
 sky130_fd_sc_hd__o21bai_1 _3936_ (.A1(_0146_),
    .A2(_0150_),
    .B1_N(_2300_),
    .Y(_0151_));
 sky130_fd_sc_hd__a21oi_2 _3937_ (.A1(_0151_),
    .A2(_2298_),
    .B1(_2297_),
    .Y(_0152_));
 sky130_fd_sc_hd__o21ai_0 _3938_ (.A1(_2295_),
    .A2(_2294_),
    .B1(_2292_),
    .Y(_0153_));
 sky130_fd_sc_hd__a31oi_4 _3939_ (.A1(_0149_),
    .A2(_0141_),
    .A3(_0152_),
    .B1(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__xnor2_1 _3940_ (.A(_0045_),
    .B(_2093_),
    .Y(_0155_));
 sky130_fd_sc_hd__o21ai_0 _3941_ (.A1(_2289_),
    .A2(_2288_),
    .B1(_2286_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21bai_1 _3942_ (.A1(_0155_),
    .A2(_0156_),
    .B1_N(_2225_),
    .Y(_0157_));
 sky130_fd_sc_hd__o41a_4 _3943_ (.A1(_2225_),
    .A2(_2288_),
    .A3(_0154_),
    .A4(_2291_),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__inv_6 _3944_ (.A(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__buf_6 _3945_ (.A(_0159_),
    .X(_2443_));
 sky130_fd_sc_hd__a21o_1 _3946_ (.A1(_2236_),
    .A2(_2331_),
    .B1(_2235_),
    .X(_0160_));
 sky130_fd_sc_hd__a21oi_1 _3947_ (.A1(_2230_),
    .A2(_0160_),
    .B1(_2229_),
    .Y(_0161_));
 sky130_fd_sc_hd__xnor2_2 _3948_ (.A(_2319_),
    .B(_0161_),
    .Y(_2320_));
 sky130_fd_sc_hd__inv_1 _3949_ (.A(_2320_),
    .Y(_2427_));
 sky130_fd_sc_hd__a21o_1 _3950_ (.A1(_2112_),
    .A2(_2333_),
    .B1(_2332_),
    .X(_0162_));
 sky130_fd_sc_hd__a21oi_2 _3951_ (.A1(_2326_),
    .A2(_0162_),
    .B1(_2325_),
    .Y(_0163_));
 sky130_fd_sc_hd__xnor2_1 _3952_ (.A(_2323_),
    .B(_0163_),
    .Y(_2336_));
 sky130_fd_sc_hd__inv_1 _3953_ (.A(_2336_),
    .Y(_2646_));
 sky130_fd_sc_hd__clkbuf_4 _3954_ (.A(_2341_),
    .X(_0164_));
 sky130_fd_sc_hd__clkinvlp_4 _3955_ (.A(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__or3_2 _3956_ (.A(_2248_),
    .B(_2240_),
    .C(_2256_),
    .X(_0166_));
 sky130_fd_sc_hd__o211ai_1 _3957_ (.A1(_0051_),
    .A2(_2248_),
    .B1(_0066_),
    .C1(_0057_),
    .Y(_0167_));
 sky130_fd_sc_hd__a21oi_1 _3958_ (.A1(_0066_),
    .A2(_2240_),
    .B1(_2256_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _3959_ (.A(_0167_),
    .B(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__o31ai_2 _3960_ (.A1(_2210_),
    .A2(_0022_),
    .A3(_0166_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__xnor2_1 _3961_ (.A(_0165_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2b_1 _3962_ (.A(_2253_),
    .B_N(_2249_),
    .Y(_0172_));
 sky130_fd_sc_hd__nor3_2 _3963_ (.A(_0046_),
    .B(_2257_),
    .C(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__nand2b_1 _3964_ (.A_N(_2245_),
    .B(_0046_),
    .Y(_0174_));
 sky130_fd_sc_hd__o311a_2 _3965_ (.A1(_2245_),
    .A2(_2253_),
    .A3(_0060_),
    .B1(_0174_),
    .C1(_0073_),
    .X(_0175_));
 sky130_fd_sc_hd__a211oi_2 _3966_ (.A1(_0055_),
    .A2(_0173_),
    .B1(_0175_),
    .C1(_2261_),
    .Y(_0176_));
 sky130_fd_sc_hd__xnor2_2 _3967_ (.A(_0165_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _3968_ (.A(_0016_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__a21oi_1 _3969_ (.A1(_0016_),
    .A2(_0171_),
    .B1(_0178_),
    .Y(_2356_));
 sky130_fd_sc_hd__clkbuf_4 _3970_ (.A(_2349_),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_1 _3971_ (.A(_2251_),
    .B(_2243_),
    .Y(_0180_));
 sky130_fd_sc_hd__a21oi_1 _3972_ (.A1(_0164_),
    .A2(_2259_),
    .B1(_2343_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_1 _3973_ (.A(_0180_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o211ai_1 _3974_ (.A1(_0057_),
    .A2(_2243_),
    .B1(_0066_),
    .C1(_0164_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _3975_ (.A(_0181_),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__o21ai_0 _3976_ (.A1(_0070_),
    .A2(_0182_),
    .B1(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__nor2b_1 _3977_ (.A(_2245_),
    .B_N(_0046_),
    .Y(_0186_));
 sky130_fd_sc_hd__o21bai_1 _3978_ (.A1(_0066_),
    .A2(_0186_),
    .B1_N(_2261_),
    .Y(_0187_));
 sky130_fd_sc_hd__a21o_1 _3979_ (.A1(_0165_),
    .A2(_0187_),
    .B1(_2345_),
    .X(_0188_));
 sky130_fd_sc_hd__nor3_1 _3980_ (.A(_2245_),
    .B(_2261_),
    .C(_2345_),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2b_1 _3981_ (.A_N(_0076_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__a21oi_1 _3982_ (.A1(_0188_),
    .A2(_0190_),
    .B1(_0009_),
    .Y(_0191_));
 sky130_fd_sc_hd__o21bai_2 _3983_ (.A1(_0013_),
    .A2(_0185_),
    .B1_N(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__xor2_4 _3984_ (.A(_0179_),
    .B(_0192_),
    .X(_2384_));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(_2213_),
    .B(_0067_),
    .Y(_0193_));
 sky130_fd_sc_hd__o21a_1 _3986_ (.A1(_0051_),
    .A2(_2251_),
    .B1(_0057_),
    .X(_0194_));
 sky130_fd_sc_hd__o21ai_0 _3987_ (.A1(_2243_),
    .A2(_0194_),
    .B1(_0066_),
    .Y(_0195_));
 sky130_fd_sc_hd__a21oi_1 _3988_ (.A1(_0095_),
    .A2(_0193_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _3989_ (.A(_2259_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__xnor2_1 _3990_ (.A(_0165_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_1 _3991_ (.A(net176),
    .B(_0177_),
    .Y(_0199_));
 sky130_fd_sc_hd__a21oi_2 _3992_ (.A1(net176),
    .A2(_0198_),
    .B1(_0199_),
    .Y(_2388_));
 sky130_fd_sc_hd__nor3_1 _3993_ (.A(_0010_),
    .B(_0078_),
    .C(_0177_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _3994_ (.A(_2213_),
    .B(_2259_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor3_1 _3995_ (.A(_2243_),
    .B(_2259_),
    .C(_0194_),
    .Y(_0202_));
 sky130_fd_sc_hd__a31oi_1 _3996_ (.A1(_0180_),
    .A2(_0095_),
    .A3(_0201_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__xnor2_1 _3997_ (.A(_0164_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__and4_1 _3998_ (.A(_0066_),
    .B(_0009_),
    .C(_0071_),
    .D(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_1 _3999_ (.A(_0164_),
    .B(_2259_),
    .X(_0206_));
 sky130_fd_sc_hd__nor4_1 _4000_ (.A(_0066_),
    .B(_0013_),
    .C(_0071_),
    .D(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__o31ai_2 _4001_ (.A1(_0200_),
    .A2(_0205_),
    .A3(_0207_),
    .B1(_0106_),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(_0115_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__xor2_1 _4003_ (.A(_2384_),
    .B(_0209_),
    .X(_2355_));
 sky130_fd_sc_hd__or2_0 _4004_ (.A(_2248_),
    .B(_0112_),
    .X(_0210_));
 sky130_fd_sc_hd__o211ai_1 _4005_ (.A1(_2248_),
    .A2(_0112_),
    .B1(_0073_),
    .C1(_0057_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor3_1 _4006_ (.A(_0057_),
    .B(_0073_),
    .C(_2240_),
    .Y(_0212_));
 sky130_fd_sc_hd__a21oi_1 _4007_ (.A1(_0073_),
    .A2(_2240_),
    .B1(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__o311a_1 _4008_ (.A1(_0073_),
    .A2(_2240_),
    .A3(_0210_),
    .B1(_0211_),
    .C1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_0016_),
    .B(_0078_),
    .Y(_0215_));
 sky130_fd_sc_hd__a21oi_1 _4010_ (.A1(_0016_),
    .A2(_0214_),
    .B1(_0215_),
    .Y(_2360_));
 sky130_fd_sc_hd__nor3_1 _4011_ (.A(_2392_),
    .B(_2396_),
    .C(_0118_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2b_1 _4012_ (.A_N(_0216_),
    .B(_0045_),
    .Y(_0217_));
 sky130_fd_sc_hd__xor2_1 _4013_ (.A(_2388_),
    .B(_0217_),
    .X(_2359_));
 sky130_fd_sc_hd__o21ai_1 _4014_ (.A1(_2265_),
    .A2(_0137_),
    .B1(_2362_),
    .Y(_0218_));
 sky130_fd_sc_hd__nor2b_1 _4015_ (.A(_2361_),
    .B_N(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__xnor2_2 _4016_ (.A(_2358_),
    .B(_0219_),
    .Y(_2404_));
 sky130_fd_sc_hd__a2111o_1 _4017_ (.A1(_2341_),
    .A2(_2256_),
    .B1(_2340_),
    .C1(_2240_),
    .D1(_2248_),
    .X(_0220_));
 sky130_fd_sc_hd__o211ai_1 _4018_ (.A1(_0046_),
    .A2(_2240_),
    .B1(_2341_),
    .C1(_0066_),
    .Y(_0221_));
 sky130_fd_sc_hd__a21oi_1 _4019_ (.A1(_2341_),
    .A2(_2256_),
    .B1(_2340_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_0221_),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__and2_1 _4021_ (.A(_2349_),
    .B(_2373_),
    .X(_0224_));
 sky130_fd_sc_hd__o211a_1 _4022_ (.A1(_0112_),
    .A2(_0220_),
    .B1(_0223_),
    .C1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__buf_4 _4023_ (.A(_2373_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _4024_ (.A1(_0226_),
    .A2(_2348_),
    .B1(_2372_),
    .X(_0227_));
 sky130_fd_sc_hd__o21ai_0 _4025_ (.A1(_0225_),
    .A2(_0227_),
    .B1(_0012_),
    .Y(_0228_));
 sky130_fd_sc_hd__buf_2 _4026_ (.A(_2377_),
    .X(_0229_));
 sky130_fd_sc_hd__nor2b_2 _4027_ (.A(_2373_),
    .B_N(_2353_),
    .Y(_0230_));
 sky130_fd_sc_hd__nor2_1 _4028_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__or3_1 _4029_ (.A(_2245_),
    .B(_2261_),
    .C(_2345_),
    .X(_0232_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(_2345_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor3b_1 _4031_ (.A(_2261_),
    .B(_2345_),
    .C_N(_2257_),
    .Y(_0234_));
 sky130_fd_sc_hd__a2111oi_4 _4032_ (.A1(_2341_),
    .A2(_0233_),
    .B1(_2349_),
    .C1(_2373_),
    .D1(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_0046_),
    .B(_0189_),
    .Y(_0236_));
 sky130_fd_sc_hd__o211ai_1 _4034_ (.A1(_0076_),
    .A2(_0232_),
    .B1(_0235_),
    .C1(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand3_1 _4035_ (.A(_0008_),
    .B(_0231_),
    .C(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__clkbuf_4 _4036_ (.A(_2365_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_1 _4037_ (.A(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21oi_1 _4038_ (.A1(_0228_),
    .A2(_0238_),
    .B1(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__and3_1 _4039_ (.A(_0240_),
    .B(_0228_),
    .C(_0238_),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_1 _4040_ (.A(_0241_),
    .B(_0242_),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2b_1 _4041_ (.A_N(_2349_),
    .B(_2345_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2b_2 _4042_ (.A_N(_2353_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__o21bai_1 _4043_ (.A1(_0164_),
    .A2(_0179_),
    .B1_N(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a2111o_1 _4044_ (.A1(_0055_),
    .A2(_0173_),
    .B1(_0175_),
    .C1(_0244_),
    .D1(_2261_),
    .X(_0246_));
 sky130_fd_sc_hd__nand3_1 _4045_ (.A(_0009_),
    .B(_0245_),
    .C(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_0164_),
    .B(_0179_),
    .Y(_0248_));
 sky130_fd_sc_hd__a21oi_1 _4047_ (.A1(_0179_),
    .A2(_2340_),
    .B1(_2348_),
    .Y(_0249_));
 sky130_fd_sc_hd__o211ai_1 _4048_ (.A1(_0170_),
    .A2(_0248_),
    .B1(_0249_),
    .C1(_0012_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand3b_1 _4049_ (.A_N(_0226_),
    .B(_0247_),
    .C(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21bo_1 _4050_ (.A1(_0247_),
    .A2(_0250_),
    .B1_N(_0226_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_0 _4051_ (.A(_0251_),
    .B(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__inv_1 _4052_ (.A(_0253_),
    .Y(_2502_));
 sky130_fd_sc_hd__a21oi_1 _4053_ (.A1(_0188_),
    .A2(_0190_),
    .B1(_0007_),
    .Y(_0254_));
 sky130_fd_sc_hd__o21ai_0 _4054_ (.A1(_0112_),
    .A2(_0220_),
    .B1(_0223_),
    .Y(_0255_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(_0008_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor3_1 _4056_ (.A(_0179_),
    .B(_0254_),
    .C(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21a_1 _4057_ (.A1(_0254_),
    .A2(_0256_),
    .B1(_0179_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _4058_ (.A(_0257_),
    .B(_0258_),
    .Y(_2506_));
 sky130_fd_sc_hd__nor2b_1 _4059_ (.A(_0181_),
    .B_N(_0179_),
    .Y(_0259_));
 sky130_fd_sc_hd__a311oi_1 _4060_ (.A1(_0164_),
    .A2(_0179_),
    .A3(_0196_),
    .B1(_0259_),
    .C1(_2351_),
    .Y(_0260_));
 sky130_fd_sc_hd__and3_1 _4061_ (.A(_0012_),
    .B(_0245_),
    .C(_0246_),
    .X(_0261_));
 sky130_fd_sc_hd__a21oi_2 _4062_ (.A1(_0009_),
    .A2(_0260_),
    .B1(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xor2_4 _4063_ (.A(_0226_),
    .B(_0262_),
    .X(_2379_));
 sky130_fd_sc_hd__inv_1 _4064_ (.A(_2382_),
    .Y(_0263_));
 sky130_fd_sc_hd__and3_1 _4065_ (.A(_2230_),
    .B(_2319_),
    .C(_0160_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(_2393_),
    .B(_2397_),
    .Y(_0265_));
 sky130_fd_sc_hd__a21oi_1 _4067_ (.A1(_2319_),
    .A2(_2229_),
    .B1(_2318_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3b_1 _4068_ (.A_N(_2401_),
    .B(_0265_),
    .C(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__buf_2 _4069_ (.A(_2402_),
    .X(_0268_));
 sky130_fd_sc_hd__o21ai_0 _4070_ (.A1(_0268_),
    .A2(_2401_),
    .B1(_2398_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor2_1 _4071_ (.A(_2394_),
    .B(_2393_),
    .Y(_0270_));
 sky130_fd_sc_hd__a21oi_1 _4072_ (.A1(_0265_),
    .A2(_0269_),
    .B1(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21ai_4 _4073_ (.A1(_0264_),
    .A2(_0267_),
    .B1(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _4074_ (.A(_2386_),
    .B(_2390_),
    .Y(_0273_));
 sky130_fd_sc_hd__a21oi_1 _4075_ (.A1(_2386_),
    .A2(_2389_),
    .B1(_2385_),
    .Y(_0274_));
 sky130_fd_sc_hd__o21ai_1 _4076_ (.A1(_0272_),
    .A2(_0273_),
    .B1(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__xnor2_2 _4077_ (.A(_0263_),
    .B(_0275_),
    .Y(_2594_));
 sky130_fd_sc_hd__nor2b_1 _4078_ (.A(_2097_),
    .B_N(_2230_),
    .Y(_0276_));
 sky130_fd_sc_hd__o2111ai_4 _4079_ (.A1(_2229_),
    .A2(_0276_),
    .B1(_2319_),
    .C1(_2398_),
    .D1(_0268_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21o_1 _4080_ (.A1(_0268_),
    .A2(_2318_),
    .B1(_2401_),
    .X(_0278_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(_2398_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__a31oi_4 _4082_ (.A1(_0265_),
    .A2(_0277_),
    .A3(_0279_),
    .B1(_0270_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_2 _4083_ (.A1(_2390_),
    .A2(_0280_),
    .B1(_2389_),
    .Y(_0281_));
 sky130_fd_sc_hd__xnor2_4 _4084_ (.A(_2386_),
    .B(_0281_),
    .Y(_2598_));
 sky130_fd_sc_hd__xnor2_2 _4085_ (.A(_2390_),
    .B(_0272_),
    .Y(_2602_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(_0277_),
    .B(_0279_),
    .Y(_0282_));
 sky130_fd_sc_hd__nor2_2 _4087_ (.A(_2397_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__xnor2_4 _4088_ (.A(_2394_),
    .B(_0283_),
    .Y(_2606_));
 sky130_fd_sc_hd__nand2b_1 _4089_ (.A_N(_0264_),
    .B(_0266_),
    .Y(_0284_));
 sky130_fd_sc_hd__a21oi_2 _4090_ (.A1(_0268_),
    .A2(_0284_),
    .B1(_2401_),
    .Y(_0285_));
 sky130_fd_sc_hd__xnor2_4 _4091_ (.A(_2398_),
    .B(_0285_),
    .Y(_2610_));
 sky130_fd_sc_hd__inv_1 _4092_ (.A(_2230_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2b_1 _4093_ (.A_N(_2318_),
    .B(_0268_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21ai_0 _4094_ (.A1(_2229_),
    .A2(_0287_),
    .B1(_2097_),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2b_1 _4095_ (.A(_0268_),
    .B_N(_2319_),
    .Y(_0289_));
 sky130_fd_sc_hd__o21ai_0 _4096_ (.A1(_2097_),
    .A2(_0289_),
    .B1(_2230_),
    .Y(_0290_));
 sky130_fd_sc_hd__o221ai_1 _4097_ (.A1(_0268_),
    .A2(_0266_),
    .B1(_0287_),
    .B2(_2319_),
    .C1(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__a211oi_2 _4098_ (.A1(_0286_),
    .A2(_0288_),
    .B1(_0291_),
    .C1(_2320_),
    .Y(_0292_));
 sky130_fd_sc_hd__nor4b_2 _4099_ (.A(_2602_),
    .B(_2606_),
    .C(_2610_),
    .D_N(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_1 _4100_ (.A(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__buf_6 _4101_ (.A(_0158_),
    .X(_0295_));
 sky130_fd_sc_hd__o21ai_0 _4102_ (.A1(_2598_),
    .A2(_0294_),
    .B1(net18),
    .Y(_0296_));
 sky130_fd_sc_hd__xor2_1 _4103_ (.A(_2594_),
    .B(_0296_),
    .X(_2403_));
 sky130_fd_sc_hd__inv_1 _4104_ (.A(_2270_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21o_1 _4105_ (.A1(_2278_),
    .A2(_2102_),
    .B1(_2277_),
    .X(_0298_));
 sky130_fd_sc_hd__a21oi_2 _4106_ (.A1(_2274_),
    .A2(_0298_),
    .B1(_2273_),
    .Y(_0299_));
 sky130_fd_sc_hd__o21bai_1 _4107_ (.A1(_0297_),
    .A2(_0299_),
    .B1_N(_2269_),
    .Y(_0300_));
 sky130_fd_sc_hd__a21oi_1 _4108_ (.A1(_2266_),
    .A2(_0300_),
    .B1(_2265_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_2 _4109_ (.A(_2362_),
    .B(_0301_),
    .Y(_2408_));
 sky130_fd_sc_hd__o21ai_0 _4110_ (.A1(_2229_),
    .A2(_0276_),
    .B1(_2319_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2b_1 _4111_ (.A_N(_2318_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__xnor2_1 _4112_ (.A(_0268_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_1 _4113_ (.A(_0304_),
    .Y(_2478_));
 sky130_fd_sc_hd__nand2_1 _4114_ (.A(_2429_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__or4_2 _4115_ (.A(_2602_),
    .B(_2606_),
    .C(_2610_),
    .D(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _4116_ (.A(net18),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__xor2_1 _4117_ (.A(_2598_),
    .B(_0307_),
    .X(_2407_));
 sky130_fd_sc_hd__nor2_1 _4118_ (.A(_2606_),
    .B(_2610_),
    .Y(_0308_));
 sky130_fd_sc_hd__a21oi_1 _4119_ (.A1(_0292_),
    .A2(_0308_),
    .B1(net2),
    .Y(_0309_));
 sky130_fd_sc_hd__xnor2_1 _4120_ (.A(_2602_),
    .B(_0309_),
    .Y(_2411_));
 sky130_fd_sc_hd__o21ai_0 _4121_ (.A1(_2610_),
    .A2(_0305_),
    .B1(_0295_),
    .Y(_0310_));
 sky130_fd_sc_hd__xor2_1 _4122_ (.A(_2606_),
    .B(_0310_),
    .X(_2415_));
 sky130_fd_sc_hd__nor2_1 _4123_ (.A(net2),
    .B(_0292_),
    .Y(_0311_));
 sky130_fd_sc_hd__xnor2_1 _4124_ (.A(_2610_),
    .B(_0311_),
    .Y(_2419_));
 sky130_fd_sc_hd__nor2_1 _4125_ (.A(_2429_),
    .B(net2),
    .Y(_0312_));
 sky130_fd_sc_hd__xnor2_1 _4126_ (.A(_2478_),
    .B(_0312_),
    .Y(_2423_));
 sky130_fd_sc_hd__nor2_1 _4127_ (.A(_0295_),
    .B(_2427_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(_2430_),
    .A2(_0295_),
    .B1(_0313_),
    .X(_2117_));
 sky130_fd_sc_hd__inv_1 _4129_ (.A(_2117_),
    .Y(_2121_));
 sky130_fd_sc_hd__inv_1 _4130_ (.A(_2425_),
    .Y(_0314_));
 sky130_fd_sc_hd__nor2b_1 _4131_ (.A(_2116_),
    .B_N(_2432_),
    .Y(_0315_));
 sky130_fd_sc_hd__o21ai_0 _4132_ (.A1(_2431_),
    .A2(_0315_),
    .B1(_2426_),
    .Y(_0316_));
 sky130_fd_sc_hd__a21boi_1 _4133_ (.A1(_0314_),
    .A2(_0316_),
    .B1_N(_2422_),
    .Y(_0317_));
 sky130_fd_sc_hd__o21a_1 _4134_ (.A1(_2421_),
    .A2(_0317_),
    .B1(_2418_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_1 _4135_ (.A(_2417_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__xnor2_2 _4136_ (.A(_2414_),
    .B(_0319_),
    .Y(_2630_));
 sky130_fd_sc_hd__nand2b_1 _4137_ (.A_N(_2119_),
    .B(_2426_),
    .Y(_0320_));
 sky130_fd_sc_hd__a21boi_0 _4138_ (.A1(_0314_),
    .A2(_0320_),
    .B1_N(_2422_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _4139_ (.A(_2421_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__xnor2_1 _4140_ (.A(_2418_),
    .B(_0322_),
    .Y(_2634_));
 sky130_fd_sc_hd__inv_1 _4141_ (.A(_2634_),
    .Y(_2493_));
 sky130_fd_sc_hd__nand2_1 _4142_ (.A(_0314_),
    .B(_0316_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(_2422_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_2 _4144_ (.A(_0317_),
    .B(_0324_),
    .Y(_2638_));
 sky130_fd_sc_hd__inv_1 _4145_ (.A(_2638_),
    .Y(_2492_));
 sky130_fd_sc_hd__o21a_1 _4146_ (.A1(_2414_),
    .A2(_2413_),
    .B1(_2410_),
    .X(_0325_));
 sky130_fd_sc_hd__nor3_1 _4147_ (.A(_2409_),
    .B(_2413_),
    .C(_2417_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2b_1 _4148_ (.A_N(_0318_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__o21ai_1 _4149_ (.A1(_2409_),
    .A2(_0325_),
    .B1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__xnor2_2 _4150_ (.A(_2406_),
    .B(_0328_),
    .Y(_2622_));
 sky130_fd_sc_hd__inv_1 _4151_ (.A(_2110_),
    .Y(_2106_));
 sky130_fd_sc_hd__inv_1 _4152_ (.A(net69),
    .Y(_2471_));
 sky130_fd_sc_hd__nand2_1 _4153_ (.A(_2473_),
    .B(_0041_),
    .Y(_0329_));
 sky130_fd_sc_hd__o21ai_2 _4154_ (.A1(_2471_),
    .A2(_0041_),
    .B1(_0329_),
    .Y(_2474_));
 sky130_fd_sc_hd__inv_1 _4155_ (.A(_2474_),
    .Y(_2123_));
 sky130_fd_sc_hd__inv_1 _4156_ (.A(_2463_),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_1 _4157_ (.A(_2468_),
    .Y(_0331_));
 sky130_fd_sc_hd__a21o_1 _4158_ (.A1(_2476_),
    .A2(net62),
    .B1(_2475_),
    .X(_0332_));
 sky130_fd_sc_hd__a21oi_4 _4159_ (.A1(_2470_),
    .A2(_0332_),
    .B1(_2469_),
    .Y(_0333_));
 sky130_fd_sc_hd__o21bai_1 _4160_ (.A1(_0333_),
    .A2(_0331_),
    .B1_N(_2467_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21oi_2 _4161_ (.A1(_0334_),
    .A2(_2466_),
    .B1(_2465_),
    .Y(_0335_));
 sky130_fd_sc_hd__o21bai_1 _4162_ (.A1(_0335_),
    .A2(_0330_),
    .B1_N(_2462_),
    .Y(_0336_));
 sky130_fd_sc_hd__a211o_1 _4163_ (.A1(_0336_),
    .A2(_2460_),
    .B1(_2459_),
    .C1(_2456_),
    .X(_0337_));
 sky130_fd_sc_hd__o211ai_2 _4164_ (.A1(_2457_),
    .A2(_2456_),
    .B1(_0337_),
    .C1(_2454_),
    .Y(_0338_));
 sky130_fd_sc_hd__nor3_1 _4165_ (.A(_2447_),
    .B(_2450_),
    .C(_2453_),
    .Y(_0339_));
 sky130_fd_sc_hd__nor3_1 _4166_ (.A(_2451_),
    .B(_2447_),
    .C(_2450_),
    .Y(_0340_));
 sky130_fd_sc_hd__nor2_1 _4167_ (.A(_2448_),
    .B(_2447_),
    .Y(_0341_));
 sky130_fd_sc_hd__a211o_4 _4168_ (.A1(_0339_),
    .A2(_0338_),
    .B1(_0340_),
    .C1(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__nand4_4 _4169_ (.A(_2435_),
    .B(_2445_),
    .C(_2438_),
    .D(_2441_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _4170_ (.A1(_2441_),
    .A2(_2444_),
    .B1(_2440_),
    .Y(_0344_));
 sky130_fd_sc_hd__nor2b_1 _4171_ (.A(_0344_),
    .B_N(_2438_),
    .Y(_0345_));
 sky130_fd_sc_hd__o21ai_0 _4172_ (.A1(_2437_),
    .A2(_0345_),
    .B1(_2435_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2b_1 _4173_ (.A_N(_2434_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__o21bai_4 _4174_ (.A1(_0343_),
    .A2(_0342_),
    .B1_N(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_6 _4175_ (.A(net174),
    .Y(_2665_));
 sky130_fd_sc_hd__inv_1 _4176_ (.A(_2323_),
    .Y(_0349_));
 sky130_fd_sc_hd__a21oi_1 _4177_ (.A1(_2326_),
    .A2(_2114_),
    .B1(_2325_),
    .Y(_0350_));
 sky130_fd_sc_hd__o21bai_1 _4178_ (.A1(_0349_),
    .A2(_0350_),
    .B1_N(_2322_),
    .Y(_0351_));
 sky130_fd_sc_hd__xor2_1 _4179_ (.A(_2480_),
    .B(_0351_),
    .X(_2481_));
 sky130_fd_sc_hd__inv_1 _4180_ (.A(_2481_),
    .Y(_2645_));
 sky130_fd_sc_hd__a21o_1 _4181_ (.A1(_2129_),
    .A2(_2491_),
    .B1(_2490_),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_2 _4182_ (.A1(_2487_),
    .A2(_0352_),
    .B1(_2486_),
    .Y(_0353_));
 sky130_fd_sc_hd__xnor2_2 _4183_ (.A(_2484_),
    .B(_0353_),
    .Y(_2499_));
 sky130_fd_sc_hd__inv_1 _4184_ (.A(_2499_),
    .Y(_2842_));
 sky130_fd_sc_hd__clkbuf_2 _4185_ (.A(_0239_),
    .X(_0354_));
 sky130_fd_sc_hd__a21o_1 _4186_ (.A1(_0226_),
    .A2(_2351_),
    .B1(_2375_),
    .X(_0355_));
 sky130_fd_sc_hd__nor4_1 _4187_ (.A(_0354_),
    .B(_0070_),
    .C(_0182_),
    .D(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__nor3_1 _4188_ (.A(_0354_),
    .B(_0224_),
    .C(_0355_),
    .Y(_0357_));
 sky130_fd_sc_hd__a21o_1 _4189_ (.A1(_0354_),
    .A2(_0355_),
    .B1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__nor3_1 _4190_ (.A(_0354_),
    .B(_0184_),
    .C(_0355_),
    .Y(_0359_));
 sky130_fd_sc_hd__o2111a_1 _4191_ (.A1(_0070_),
    .A2(_0182_),
    .B1(_0224_),
    .C1(_0184_),
    .D1(_0354_),
    .X(_0360_));
 sky130_fd_sc_hd__or4_2 _4192_ (.A(_0356_),
    .B(_0358_),
    .C(_0359_),
    .D(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__and3_1 _4193_ (.A(_0354_),
    .B(_0235_),
    .C(_0236_),
    .X(_0362_));
 sky130_fd_sc_hd__a2111oi_2 _4194_ (.A1(_0235_),
    .A2(_0236_),
    .B1(_0354_),
    .C1(_0229_),
    .D1(_0230_),
    .Y(_0363_));
 sky130_fd_sc_hd__or3_1 _4195_ (.A(_0239_),
    .B(_0229_),
    .C(_0230_),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_0 _4196_ (.A1(_0229_),
    .A2(_0230_),
    .B1(_0354_),
    .Y(_0365_));
 sky130_fd_sc_hd__o31ai_2 _4197_ (.A1(_0076_),
    .A2(_0232_),
    .A3(_0364_),
    .B1(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a2111oi_4 _4198_ (.A1(_0190_),
    .A2(_0362_),
    .B1(_0363_),
    .C1(_0366_),
    .D1(net171),
    .Y(_0367_));
 sky130_fd_sc_hd__a21oi_2 _4199_ (.A1(net176),
    .A2(_0361_),
    .B1(_0367_),
    .Y(_2530_));
 sky130_fd_sc_hd__or3_1 _4200_ (.A(_2384_),
    .B(_0208_),
    .C(_2379_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_1 _4201_ (.A(_0115_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__xor2_1 _4202_ (.A(_2530_),
    .B(_0369_),
    .X(_2501_));
 sky130_fd_sc_hd__nor2_1 _4203_ (.A(_2384_),
    .B(_2388_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(_0216_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(_0115_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__xor2_1 _4206_ (.A(_2379_),
    .B(_0372_),
    .X(_2505_));
 sky130_fd_sc_hd__inv_1 _4207_ (.A(_2504_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _4208_ (.A(_2358_),
    .B(_2508_),
    .Y(_0374_));
 sky130_fd_sc_hd__a21o_1 _4209_ (.A1(_2358_),
    .A2(_2361_),
    .B1(_2357_),
    .X(_0375_));
 sky130_fd_sc_hd__a21oi_1 _4210_ (.A1(_2508_),
    .A2(_0375_),
    .B1(_2507_),
    .Y(_0376_));
 sky130_fd_sc_hd__o21ai_1 _4211_ (.A1(_0218_),
    .A2(_0374_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__xnor2_2 _4212_ (.A(_0373_),
    .B(_0377_),
    .Y(_2534_));
 sky130_fd_sc_hd__nor2b_1 _4213_ (.A(_2519_),
    .B_N(_2369_),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _4214_ (.A(_2523_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__a211o_1 _4215_ (.A1(_0231_),
    .A2(_0237_),
    .B1(_0239_),
    .C1(_2519_),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _4216_ (.A(_0379_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_4 _4217_ (.A(_2511_),
    .X(_0382_));
 sky130_fd_sc_hd__clkinvlp_4 _4218_ (.A(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_1 _4219_ (.A(_0383_),
    .B(_0007_),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_1 _4220_ (.A(_0382_),
    .B(_0007_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21boi_1 _4221_ (.A1(_0379_),
    .A2(_0380_),
    .B1_N(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__buf_4 _4222_ (.A(_2519_),
    .X(_0387_));
 sky130_fd_sc_hd__a21oi_1 _4223_ (.A1(_0387_),
    .A2(_2364_),
    .B1(_2518_),
    .Y(_0388_));
 sky130_fd_sc_hd__and2_0 _4224_ (.A(_0239_),
    .B(_2519_),
    .X(_0389_));
 sky130_fd_sc_hd__o21ai_0 _4225_ (.A1(_0225_),
    .A2(_0227_),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__and4_1 _4226_ (.A(_0383_),
    .B(_0007_),
    .C(_0388_),
    .D(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_0382_),
    .B(_0007_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21oi_1 _4228_ (.A1(_0388_),
    .A2(_0390_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__a2111oi_4 _4229_ (.A1(_0381_),
    .A2(_0384_),
    .B1(_0386_),
    .C1(_0391_),
    .D1(_0393_),
    .Y(_2566_));
 sky130_fd_sc_hd__nor3_1 _4230_ (.A(_2261_),
    .B(_2369_),
    .C(_0229_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand3b_1 _4231_ (.A_N(_2353_),
    .B(_0243_),
    .C(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a211oi_4 _4232_ (.A1(_0055_),
    .A2(_0173_),
    .B1(_0175_),
    .C1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_1 _4233_ (.A(_0229_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_1 _4234_ (.A1(_0226_),
    .A2(_0397_),
    .B1(_0239_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(_2369_),
    .B(_0229_),
    .Y(_0399_));
 sky130_fd_sc_hd__o21ai_1 _4236_ (.A1(_0164_),
    .A2(_2349_),
    .B1(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o22ai_4 _4237_ (.A1(_2369_),
    .A2(_0398_),
    .B1(_0400_),
    .B2(_0244_),
    .Y(_0401_));
 sky130_fd_sc_hd__or2_0 _4238_ (.A(_0396_),
    .B(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and4_1 _4239_ (.A(_0164_),
    .B(_0179_),
    .C(_0226_),
    .D(_0239_),
    .X(_0403_));
 sky130_fd_sc_hd__o311ai_4 _4240_ (.A1(_2210_),
    .A2(_0022_),
    .A3(_0166_),
    .B1(_0403_),
    .C1(_0169_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_0226_),
    .B(_0239_),
    .Y(_0405_));
 sky130_fd_sc_hd__nor2_1 _4242_ (.A(_0249_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__a211oi_2 _4243_ (.A1(_0239_),
    .A2(_2372_),
    .B1(_2364_),
    .C1(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand3_1 _4244_ (.A(_0007_),
    .B(_0404_),
    .C(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__o21ai_1 _4245_ (.A1(_0012_),
    .A2(_0402_),
    .B1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_2 _4246_ (.A(_0387_),
    .B(_0409_),
    .Y(_2574_));
 sky130_fd_sc_hd__nor2_1 _4247_ (.A(_0396_),
    .B(_0401_),
    .Y(_0410_));
 sky130_fd_sc_hd__a211o_1 _4248_ (.A1(_2343_),
    .A2(_0179_),
    .B1(_2351_),
    .C1(_2375_),
    .X(_0411_));
 sky130_fd_sc_hd__o211ai_1 _4249_ (.A1(_0226_),
    .A2(_2375_),
    .B1(_0411_),
    .C1(_0354_),
    .Y(_0412_));
 sky130_fd_sc_hd__a21oi_1 _4250_ (.A1(_2259_),
    .A2(_0403_),
    .B1(_2367_),
    .Y(_0413_));
 sky130_fd_sc_hd__nand2_1 _4251_ (.A(_0412_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__o211ai_1 _4252_ (.A1(_2243_),
    .A2(_0194_),
    .B1(_0403_),
    .C1(_0066_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21oi_2 _4253_ (.A1(_0095_),
    .A2(_0193_),
    .B1(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__or2_0 _4254_ (.A(_0414_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _4255_ (.A(_0014_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__a21oi_1 _4256_ (.A1(_0014_),
    .A2(_0410_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__xnor2_2 _4257_ (.A(_0387_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_1 _4258_ (.A(_0420_),
    .Y(_2525_));
 sky130_fd_sc_hd__nand3_1 _4259_ (.A(_2386_),
    .B(_2382_),
    .C(_2390_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21bai_1 _4260_ (.A1(_0263_),
    .A2(_0274_),
    .B1_N(_2381_),
    .Y(_0422_));
 sky130_fd_sc_hd__o21bai_1 _4261_ (.A1(_0272_),
    .A2(_0421_),
    .B1_N(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a21oi_1 _4262_ (.A1(_2532_),
    .A2(_0423_),
    .B1(_2531_),
    .Y(_0424_));
 sky130_fd_sc_hd__xnor2_2 _4263_ (.A(_2528_),
    .B(_0424_),
    .Y(_2586_));
 sky130_fd_sc_hd__a41oi_4 _4264_ (.A1(_2386_),
    .A2(_2382_),
    .A3(_2390_),
    .A4(_0280_),
    .B1(_0422_),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_2 _4265_ (.A(_2532_),
    .B(_0425_),
    .Y(_2590_));
 sky130_fd_sc_hd__nor3_1 _4266_ (.A(_2594_),
    .B(_2598_),
    .C(_2590_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21oi_1 _4267_ (.A1(_0293_),
    .A2(_0426_),
    .B1(net2),
    .Y(_0427_));
 sky130_fd_sc_hd__xnor2_1 _4268_ (.A(_2586_),
    .B(_0427_),
    .Y(_2533_));
 sky130_fd_sc_hd__a2111oi_2 _4269_ (.A1(_2266_),
    .A2(_0300_),
    .B1(_2361_),
    .C1(_2357_),
    .D1(_2265_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor3_1 _4270_ (.A(_2362_),
    .B(_2357_),
    .C(_2361_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_1 _4271_ (.A(_2358_),
    .B(_2357_),
    .Y(_0430_));
 sky130_fd_sc_hd__nor3_2 _4272_ (.A(_0428_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__xor2_4 _4273_ (.A(_2508_),
    .B(_0431_),
    .X(_2538_));
 sky130_fd_sc_hd__o31ai_1 _4274_ (.A1(_2594_),
    .A2(_2598_),
    .A3(_0306_),
    .B1(net18),
    .Y(_0432_));
 sky130_fd_sc_hd__xor2_1 _4275_ (.A(_2590_),
    .B(_0432_),
    .X(_2537_));
 sky130_fd_sc_hd__nor2_1 _4276_ (.A(_2405_),
    .B(_2539_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(_0326_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__o21ai_1 _4278_ (.A1(_2409_),
    .A2(_0325_),
    .B1(_2406_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _4279_ (.A(_0435_),
    .B(_0433_),
    .Y(_0436_));
 sky130_fd_sc_hd__o221ai_4 _4280_ (.A1(_2540_),
    .A2(_2539_),
    .B1(_0318_),
    .B2(_0434_),
    .C1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__xor2_2 _4281_ (.A(_2536_),
    .B(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__inv_1 _4282_ (.A(_0438_),
    .Y(_2614_));
 sky130_fd_sc_hd__clkbuf_4 _4283_ (.A(_2543_),
    .X(_0439_));
 sky130_fd_sc_hd__and4_1 _4284_ (.A(_0382_),
    .B(_2551_),
    .C(_0224_),
    .D(_0389_),
    .X(_0440_));
 sky130_fd_sc_hd__o211a_1 _4285_ (.A1(_0112_),
    .A2(_0220_),
    .B1(_0223_),
    .C1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_0382_),
    .B(_2551_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _4287_ (.A1(_2551_),
    .A2(_2510_),
    .B1(_2550_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_1 _4288_ (.A(_0387_),
    .Y(_0444_));
 sky130_fd_sc_hd__nor3_1 _4289_ (.A(_0240_),
    .B(_0444_),
    .C(_0442_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(_0227_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__o211ai_1 _4291_ (.A1(_0388_),
    .A2(_0442_),
    .B1(_0443_),
    .C1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor4_2 _4292_ (.A(_0239_),
    .B(_0387_),
    .C(_2511_),
    .D(_2551_),
    .Y(_0448_));
 sky130_fd_sc_hd__o2111a_1 _4293_ (.A1(_0076_),
    .A2(_0232_),
    .B1(_0235_),
    .C1(_0236_),
    .D1(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__clkinv_4 _4294_ (.A(_2551_),
    .Y(_0450_));
 sky130_fd_sc_hd__o211ai_1 _4295_ (.A1(_2523_),
    .A2(_0378_),
    .B1(_0383_),
    .C1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__a21oi_1 _4296_ (.A1(_2515_),
    .A2(_0450_),
    .B1(_2555_),
    .Y(_0452_));
 sky130_fd_sc_hd__o21ai_0 _4297_ (.A1(_0229_),
    .A2(_0230_),
    .B1(_0448_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand3_1 _4298_ (.A(_0451_),
    .B(_0452_),
    .C(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21ai_0 _4299_ (.A1(_0449_),
    .A2(_0454_),
    .B1(_0008_),
    .Y(_0455_));
 sky130_fd_sc_hd__o31ai_2 _4300_ (.A1(_0008_),
    .A2(_0441_),
    .A3(_0447_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__xnor2_2 _4301_ (.A(_0439_),
    .B(_0456_),
    .Y(_2558_));
 sky130_fd_sc_hd__o21ai_0 _4302_ (.A1(_0449_),
    .A2(_0454_),
    .B1(_0013_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand3_1 _4303_ (.A(_0387_),
    .B(_0382_),
    .C(_2367_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_2 _4304_ (.A1(_0382_),
    .A2(_2521_),
    .B1(_2513_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _4305_ (.A1(_0458_),
    .A2(_0459_),
    .B1(_0450_),
    .Y(_0460_));
 sky130_fd_sc_hd__a211oi_1 _4306_ (.A1(_0355_),
    .A2(_0445_),
    .B1(_0460_),
    .C1(_2553_),
    .Y(_0461_));
 sky130_fd_sc_hd__o211ai_1 _4307_ (.A1(_0070_),
    .A2(_0182_),
    .B1(_0440_),
    .C1(_0184_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand3_1 _4308_ (.A(net171),
    .B(_0461_),
    .C(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(_0457_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__xnor2_2 _4310_ (.A(_0439_),
    .B(_0464_),
    .Y(_2736_));
 sky130_fd_sc_hd__a21oi_1 _4311_ (.A1(_0383_),
    .A2(_2523_),
    .B1(_2515_),
    .Y(_0465_));
 sky130_fd_sc_hd__o41ai_4 _4312_ (.A1(_0387_),
    .A2(_2511_),
    .A3(_0396_),
    .A4(_0401_),
    .B1(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand3_1 _4313_ (.A(_0412_),
    .B(_0413_),
    .C(_0459_),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_0 _4314_ (.A1(_0444_),
    .A2(_0383_),
    .B1(_0459_),
    .Y(_0468_));
 sky130_fd_sc_hd__o211ai_1 _4315_ (.A1(_0416_),
    .A2(_0467_),
    .B1(_0468_),
    .C1(net171),
    .Y(_0469_));
 sky130_fd_sc_hd__o21ai_2 _4316_ (.A1(net171),
    .A2(_0466_),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__xnor2_4 _4317_ (.A(_0450_),
    .B(_0470_),
    .Y(_2724_));
 sky130_fd_sc_hd__o211ai_1 _4318_ (.A1(_0070_),
    .A2(_0182_),
    .B1(_0224_),
    .C1(_0184_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor3_1 _4319_ (.A(_2367_),
    .B(_2521_),
    .C(_0355_),
    .Y(_0472_));
 sky130_fd_sc_hd__or2_0 _4320_ (.A(_0354_),
    .B(_2367_),
    .X(_0473_));
 sky130_fd_sc_hd__a21oi_1 _4321_ (.A1(_0387_),
    .A2(_0473_),
    .B1(_2521_),
    .Y(_0474_));
 sky130_fd_sc_hd__a21oi_1 _4322_ (.A1(_0471_),
    .A2(_0472_),
    .B1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__mux2i_2 _4323_ (.A0(_0384_),
    .A1(_0385_),
    .S(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand4_1 _4324_ (.A(_0383_),
    .B(_0013_),
    .C(_0379_),
    .D(_0380_),
    .Y(_0477_));
 sky130_fd_sc_hd__o211ai_4 _4325_ (.A1(_0381_),
    .A2(_0392_),
    .B1(_0476_),
    .C1(_0477_),
    .Y(_2578_));
 sky130_fd_sc_hd__xnor2_4 _4326_ (.A(net36),
    .B(net52),
    .Y(_0478_));
 sky130_fd_sc_hd__a211oi_1 _4327_ (.A1(_0450_),
    .A2(_0466_),
    .B1(_2555_),
    .C1(_2547_),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2b_1 _4328_ (.A(_2547_),
    .B_N(_0439_),
    .Y(_0480_));
 sky130_fd_sc_hd__nor2_1 _4329_ (.A(_0414_),
    .B(_0416_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand4_1 _4330_ (.A(_0387_),
    .B(_0382_),
    .C(_2551_),
    .D(_0439_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21bai_1 _4331_ (.A1(_0450_),
    .A2(_0459_),
    .B1_N(_2553_),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_1 _4332_ (.A1(_0439_),
    .A2(_0483_),
    .B1(_2545_),
    .Y(_0484_));
 sky130_fd_sc_hd__o211ai_1 _4333_ (.A1(_0481_),
    .A2(_0482_),
    .B1(_0484_),
    .C1(net171),
    .Y(_0485_));
 sky130_fd_sc_hd__o31a_2 _4334_ (.A1(_0008_),
    .A2(_0479_),
    .A3(_0480_),
    .B1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__xnor2_1 _4335_ (.A(_0478_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor4_1 _4336_ (.A(_2379_),
    .B(_2530_),
    .C(_0371_),
    .D(_2578_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_0420_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o31ai_1 _4338_ (.A1(_2736_),
    .A2(_2724_),
    .A3(_0489_),
    .B1(_0115_),
    .Y(_0490_));
 sky130_fd_sc_hd__xnor2_1 _4339_ (.A(_0487_),
    .B(_0490_),
    .Y(_2557_));
 sky130_fd_sc_hd__a21oi_1 _4340_ (.A1(_0382_),
    .A2(_2518_),
    .B1(_2510_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_0 _4341_ (.A1(_0387_),
    .A2(_2518_),
    .B1(_0382_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_1 _4342_ (.A(_2510_),
    .Y(_0493_));
 sky130_fd_sc_hd__a32o_1 _4343_ (.A1(_0404_),
    .A2(_0407_),
    .A3(_0491_),
    .B1(_0492_),
    .B2(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2i_2 _4344_ (.A0(_0466_),
    .A1(_0494_),
    .S(_0012_),
    .Y(_0495_));
 sky130_fd_sc_hd__xnor2_2 _4345_ (.A(_0450_),
    .B(_0495_),
    .Y(_2562_));
 sky130_fd_sc_hd__nor3_1 _4346_ (.A(_2384_),
    .B(_0208_),
    .C(_2379_),
    .Y(_0496_));
 sky130_fd_sc_hd__a32oi_1 _4347_ (.A1(net176),
    .A2(_0361_),
    .A3(_0417_),
    .B1(_0402_),
    .B2(_0367_),
    .Y(_0497_));
 sky130_fd_sc_hd__a32oi_1 _4348_ (.A1(net176),
    .A2(_0361_),
    .A3(_0481_),
    .B1(_0410_),
    .B2(_0367_),
    .Y(_0498_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(_0497_),
    .A1(_0498_),
    .S(_0444_),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_1 _4350_ (.A(_2578_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _4351_ (.A(_0496_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__o21ai_1 _4352_ (.A1(_2724_),
    .A2(_0501_),
    .B1(net4),
    .Y(_0502_));
 sky130_fd_sc_hd__xor2_1 _4353_ (.A(_2736_),
    .B(_0502_),
    .X(_2561_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_0115_),
    .B(_0489_),
    .Y(_0503_));
 sky130_fd_sc_hd__xor2_1 _4355_ (.A(_2724_),
    .B(_0503_),
    .X(_2565_));
 sky130_fd_sc_hd__o21ai_0 _4356_ (.A1(_0368_),
    .A2(_0499_),
    .B1(net4),
    .Y(_0504_));
 sky130_fd_sc_hd__xor2_1 _4357_ (.A(_2578_),
    .B(_0504_),
    .X(_2573_));
 sky130_fd_sc_hd__o31ai_1 _4358_ (.A1(_2379_),
    .A2(_2530_),
    .A3(_0371_),
    .B1(_0125_),
    .Y(_0505_));
 sky130_fd_sc_hd__xnor2_1 _4359_ (.A(_0420_),
    .B(_0505_),
    .Y(_2569_));
 sky130_fd_sc_hd__a21o_1 _4360_ (.A1(_2508_),
    .A2(_2357_),
    .B1(_2507_),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _4361_ (.A1(_2504_),
    .A2(_0506_),
    .B1(_2503_),
    .Y(_0507_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(_2265_),
    .B(_2361_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _4363_ (.A(_0507_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__a21oi_1 _4364_ (.A1(_2266_),
    .A2(_0300_),
    .B1(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nor2_1 _4365_ (.A(_2362_),
    .B(_2361_),
    .Y(_0511_));
 sky130_fd_sc_hd__o31a_1 _4366_ (.A1(_0373_),
    .A2(_0374_),
    .A3(_0511_),
    .B1(_0507_),
    .X(_0512_));
 sky130_fd_sc_hd__nand3_1 _4367_ (.A(_2576_),
    .B(_2568_),
    .C(_2572_),
    .Y(_0513_));
 sky130_fd_sc_hd__nor3_1 _4368_ (.A(_0510_),
    .B(_0512_),
    .C(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__and3_1 _4369_ (.A(_2576_),
    .B(_2568_),
    .C(_2571_),
    .X(_0515_));
 sky130_fd_sc_hd__a2111o_1 _4370_ (.A1(_2568_),
    .A2(_2575_),
    .B1(_0514_),
    .C1(_0515_),
    .D1(_2567_),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_1 _4371_ (.A1(_2564_),
    .A2(_0516_),
    .B1(_2563_),
    .Y(_0517_));
 sky130_fd_sc_hd__xnor2_2 _4372_ (.A(_2560_),
    .B(_0517_),
    .Y(_2756_));
 sky130_fd_sc_hd__nor2_1 _4373_ (.A(_0373_),
    .B(_0374_),
    .Y(_0518_));
 sky130_fd_sc_hd__o211ai_1 _4374_ (.A1(_2265_),
    .A2(_0137_),
    .B1(_0518_),
    .C1(_2362_),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_1 _4375_ (.A(_0373_),
    .B(_0376_),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(_2503_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__clkinvlp_4 _4377_ (.A(_2572_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21o_1 _4378_ (.A1(_0519_),
    .A2(_0521_),
    .B1(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__nor2_1 _4379_ (.A(_2571_),
    .B(_2575_),
    .Y(_0524_));
 sky130_fd_sc_hd__o21ai_0 _4380_ (.A1(_2576_),
    .A2(_2575_),
    .B1(_2568_),
    .Y(_0525_));
 sky130_fd_sc_hd__a21oi_1 _4381_ (.A1(_0523_),
    .A2(_0524_),
    .B1(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__or2_1 _4382_ (.A(_2567_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__xor2_2 _4383_ (.A(_2564_),
    .B(_0527_),
    .X(_2764_));
 sky130_fd_sc_hd__inv_1 _4384_ (.A(_2571_),
    .Y(_0528_));
 sky130_fd_sc_hd__o31ai_1 _4385_ (.A1(_0522_),
    .A2(_0510_),
    .A3(_0512_),
    .B1(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21oi_1 _4386_ (.A1(_2576_),
    .A2(_0529_),
    .B1(_2575_),
    .Y(_0530_));
 sky130_fd_sc_hd__xnor2_2 _4387_ (.A(_2568_),
    .B(_0530_),
    .Y(_2760_));
 sky130_fd_sc_hd__nand2_1 _4388_ (.A(_0528_),
    .B(_0523_),
    .Y(_0531_));
 sky130_fd_sc_hd__xor2_4 _4389_ (.A(_2576_),
    .B(_0531_),
    .X(_2728_));
 sky130_fd_sc_hd__nor2_1 _4390_ (.A(_0510_),
    .B(_0512_),
    .Y(_0532_));
 sky130_fd_sc_hd__xnor2_4 _4391_ (.A(_0522_),
    .B(_0532_),
    .Y(_2732_));
 sky130_fd_sc_hd__o21ai_1 _4392_ (.A1(_2532_),
    .A2(_2531_),
    .B1(_2528_),
    .Y(_0533_));
 sky130_fd_sc_hd__nor2b_1 _4393_ (.A(_2531_),
    .B_N(_0425_),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_1 _4394_ (.A(_2527_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_1 _4395_ (.A1(_0533_),
    .A2(_0534_),
    .B1(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__xnor2_2 _4396_ (.A(_2580_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_1 _4397_ (.A(_0537_),
    .Y(_2581_));
 sky130_fd_sc_hd__a21oi_2 _4398_ (.A1(_2480_),
    .A2(_0351_),
    .B1(_2479_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand3_1 _4399_ (.A(_2604_),
    .B(_2608_),
    .C(_2612_),
    .Y(_0539_));
 sky130_fd_sc_hd__a21o_1 _4400_ (.A1(_2604_),
    .A2(_2607_),
    .B1(_2603_),
    .X(_0540_));
 sky130_fd_sc_hd__a31oi_2 _4401_ (.A1(_2604_),
    .A2(_2608_),
    .A3(_2611_),
    .B1(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__o21ai_4 _4402_ (.A1(_0538_),
    .A2(_0539_),
    .B1(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand3_1 _4403_ (.A(_2592_),
    .B(_2596_),
    .C(_2599_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_2592_),
    .B(_2595_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a41oi_4 _4406_ (.A1(_2592_),
    .A2(_2596_),
    .A3(_2600_),
    .A4(_0542_),
    .B1(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nor3_1 _4407_ (.A(_2584_),
    .B(_2587_),
    .C(_2591_),
    .Y(_0547_));
 sky130_fd_sc_hd__nor3_1 _4408_ (.A(_2584_),
    .B(_2588_),
    .C(_2587_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _4409_ (.A(_2587_),
    .B(_2591_),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_1 _4410_ (.A1(_2588_),
    .A2(_2587_),
    .B1(_2584_),
    .Y(_0550_));
 sky130_fd_sc_hd__a21oi_2 _4411_ (.A1(_0546_),
    .A2(_0549_),
    .B1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__a211oi_4 _4412_ (.A1(_0546_),
    .A2(_0547_),
    .B1(_0548_),
    .C1(_0551_),
    .Y(_2772_));
 sky130_fd_sc_hd__nor2_1 _4413_ (.A(_2595_),
    .B(_2599_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor3_1 _4414_ (.A(_2322_),
    .B(_2479_),
    .C(_2611_),
    .Y(_0553_));
 sky130_fd_sc_hd__o21ai_1 _4415_ (.A1(_0349_),
    .A2(_0163_),
    .B1(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_1 _4416_ (.A(_2612_),
    .Y(_0555_));
 sky130_fd_sc_hd__nor2_1 _4417_ (.A(_2480_),
    .B(_2479_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_1 _4418_ (.A(_2611_),
    .Y(_0557_));
 sky130_fd_sc_hd__o21ai_1 _4419_ (.A1(_0555_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__a41oi_2 _4420_ (.A1(_2604_),
    .A2(_2608_),
    .A3(_0554_),
    .A4(_0558_),
    .B1(_0540_),
    .Y(_0559_));
 sky130_fd_sc_hd__o21a_1 _4421_ (.A1(_2600_),
    .A2(_2599_),
    .B1(_2596_),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_1 _4422_ (.A(_2595_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _4423_ (.A1(_0552_),
    .A2(_0559_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a21oi_1 _4424_ (.A1(_2592_),
    .A2(_0562_),
    .B1(_2591_),
    .Y(_0563_));
 sky130_fd_sc_hd__xnor2_2 _4425_ (.A(_2588_),
    .B(_0563_),
    .Y(_2802_));
 sky130_fd_sc_hd__a21o_1 _4426_ (.A1(_2600_),
    .A2(_0542_),
    .B1(_2599_),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _4427_ (.A1(_2596_),
    .A2(_0564_),
    .B1(_2595_),
    .Y(_0565_));
 sky130_fd_sc_hd__xnor2_2 _4428_ (.A(_2592_),
    .B(_0565_),
    .Y(_2778_));
 sky130_fd_sc_hd__nor2b_1 _4429_ (.A(_0559_),
    .B_N(_2600_),
    .Y(_0566_));
 sky130_fd_sc_hd__nor2_1 _4430_ (.A(_2599_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__xnor2_2 _4431_ (.A(_2596_),
    .B(_0567_),
    .Y(_2782_));
 sky130_fd_sc_hd__xor2_2 _4432_ (.A(_2600_),
    .B(_0542_),
    .X(_2786_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(_2646_),
    .B(_2645_),
    .Y(_0568_));
 sky130_fd_sc_hd__a31oi_2 _4434_ (.A1(_2608_),
    .A2(_0554_),
    .A3(_0558_),
    .B1(_2607_),
    .Y(_0569_));
 sky130_fd_sc_hd__xnor2_2 _4435_ (.A(_2604_),
    .B(_0569_),
    .Y(_2790_));
 sky130_fd_sc_hd__o21ai_1 _4436_ (.A1(_0555_),
    .A2(_0538_),
    .B1(_0557_),
    .Y(_0570_));
 sky130_fd_sc_hd__xnor2_2 _4437_ (.A(_2608_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__o21bai_1 _4438_ (.A1(_0349_),
    .A2(_0163_),
    .B1_N(_2322_),
    .Y(_0572_));
 sky130_fd_sc_hd__a21oi_1 _4439_ (.A1(_2480_),
    .A2(_0572_),
    .B1(_2479_),
    .Y(_0573_));
 sky130_fd_sc_hd__xnor2_1 _4440_ (.A(_0555_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_0571_),
    .B(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__nor3_1 _4442_ (.A(_2786_),
    .B(_2790_),
    .C(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__or4b_1 _4443_ (.A(_2802_),
    .B(_2778_),
    .C(_2782_),
    .D_N(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__buf_2 _4444_ (.A(net174),
    .X(_0578_));
 sky130_fd_sc_hd__o21ai_0 _4445_ (.A1(_0568_),
    .A2(_0577_),
    .B1(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__xor2_1 _4446_ (.A(_2772_),
    .B(_0579_),
    .X(_2613_));
 sky130_fd_sc_hd__inv_1 _4447_ (.A(_0574_),
    .Y(_2696_));
 sky130_fd_sc_hd__inv_1 _4448_ (.A(_2647_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2b_1 _4449_ (.A_N(_2782_),
    .B(_0576_),
    .Y(_0581_));
 sky130_fd_sc_hd__o31a_1 _4450_ (.A1(_0580_),
    .A2(_2778_),
    .A3(_0581_),
    .B1(net6),
    .X(_0582_));
 sky130_fd_sc_hd__xnor2_1 _4451_ (.A(_2802_),
    .B(_0582_),
    .Y(_2617_));
 sky130_fd_sc_hd__o21ai_0 _4452_ (.A1(_0568_),
    .A2(_0581_),
    .B1(_0578_),
    .Y(_0583_));
 sky130_fd_sc_hd__xor2_1 _4453_ (.A(_2778_),
    .B(_0583_),
    .X(_2621_));
 sky130_fd_sc_hd__a21oi_1 _4454_ (.A1(_2647_),
    .A2(_0576_),
    .B1(_2665_),
    .Y(_0584_));
 sky130_fd_sc_hd__xnor2_1 _4455_ (.A(_2782_),
    .B(_0584_),
    .Y(_2625_));
 sky130_fd_sc_hd__o31ai_1 _4456_ (.A1(_0568_),
    .A2(_2790_),
    .A3(_0575_),
    .B1(_0578_),
    .Y(_0585_));
 sky130_fd_sc_hd__xor2_1 _4457_ (.A(_2786_),
    .B(_0585_),
    .X(_2629_));
 sky130_fd_sc_hd__o21ai_0 _4458_ (.A1(_0580_),
    .A2(_0575_),
    .B1(net174),
    .Y(_0586_));
 sky130_fd_sc_hd__xor2_1 _4459_ (.A(_2790_),
    .B(_0586_),
    .X(_2633_));
 sky130_fd_sc_hd__o21ai_0 _4460_ (.A1(_0568_),
    .A2(_2696_),
    .B1(_0578_),
    .Y(_0587_));
 sky130_fd_sc_hd__xnor2_1 _4461_ (.A(_0571_),
    .B(_0587_),
    .Y(_2637_));
 sky130_fd_sc_hd__nor2_1 _4462_ (.A(_2647_),
    .B(_2665_),
    .Y(_0588_));
 sky130_fd_sc_hd__xnor2_1 _4463_ (.A(_2696_),
    .B(_0588_),
    .Y(_2641_));
 sky130_fd_sc_hd__buf_6 _4464_ (.A(_0348_),
    .X(_2652_));
 sky130_fd_sc_hd__nor2_1 _4465_ (.A(net9),
    .B(_2645_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_2 _4466_ (.A1(_2648_),
    .A2(net9),
    .B1(_0589_),
    .Y(_2132_));
 sky130_fd_sc_hd__inv_1 _4467_ (.A(_2627_),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_1 _4468_ (.A(_2635_),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_1 _4469_ (.A(_2643_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2b_1 _4470_ (.A(_2337_),
    .B_N(_2650_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_0 _4471_ (.A1(_2649_),
    .A2(_0593_),
    .B1(_2644_),
    .Y(_0594_));
 sky130_fd_sc_hd__a21boi_0 _4472_ (.A1(_0592_),
    .A2(_0594_),
    .B1_N(_2640_),
    .Y(_0595_));
 sky130_fd_sc_hd__o21ai_0 _4473_ (.A1(_2639_),
    .A2(_0595_),
    .B1(_2636_),
    .Y(_0596_));
 sky130_fd_sc_hd__a21boi_0 _4474_ (.A1(_0591_),
    .A2(_0596_),
    .B1_N(_2632_),
    .Y(_0597_));
 sky130_fd_sc_hd__o21ai_1 _4475_ (.A1(_2631_),
    .A2(_0597_),
    .B1(_2628_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3_1 _4476_ (.A(_2624_),
    .B(_2620_),
    .C(_2616_),
    .Y(_0599_));
 sky130_fd_sc_hd__a21o_1 _4477_ (.A1(_0590_),
    .A2(_0598_),
    .B1(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__and3_1 _4478_ (.A(_2620_),
    .B(_2616_),
    .C(_2623_),
    .X(_0601_));
 sky130_fd_sc_hd__a21oi_1 _4479_ (.A1(_2616_),
    .A2(_2619_),
    .B1(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_0600_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_2 _4481_ (.A(_0590_),
    .B(_0598_),
    .Y(_0604_));
 sky130_fd_sc_hd__a21o_1 _4482_ (.A1(_2624_),
    .A2(_0604_),
    .B1(_2623_),
    .X(_0605_));
 sky130_fd_sc_hd__a211oi_1 _4483_ (.A1(_2620_),
    .A2(_0605_),
    .B1(_2619_),
    .C1(_2616_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_2 _4484_ (.A(_0603_),
    .B(_0606_),
    .Y(_2848_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(_0591_),
    .B(_0596_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_1 _4486_ (.A(_2632_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_1 _4487_ (.A(_0597_),
    .B(_0608_),
    .Y(_2826_));
 sky130_fd_sc_hd__inv_1 _4488_ (.A(_2826_),
    .Y(_2715_));
 sky130_fd_sc_hd__a21o_1 _4489_ (.A1(_2134_),
    .A2(_2644_),
    .B1(_2643_),
    .X(_0609_));
 sky130_fd_sc_hd__a21oi_1 _4490_ (.A1(_2640_),
    .A2(_0609_),
    .B1(_2639_),
    .Y(_0610_));
 sky130_fd_sc_hd__xnor2_2 _4491_ (.A(_2636_),
    .B(_0610_),
    .Y(_2830_));
 sky130_fd_sc_hd__inv_1 _4492_ (.A(_2830_),
    .Y(_2714_));
 sky130_fd_sc_hd__inv_1 _4493_ (.A(_2678_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_1 _4494_ (.A(_2684_),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_1 _4495_ (.A(_2690_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2b_1 _4496_ (.A(net62),
    .B_N(_2694_),
    .Y(_0614_));
 sky130_fd_sc_hd__o21ai_1 _4497_ (.A1(_0614_),
    .A2(_2693_),
    .B1(_2691_),
    .Y(_0615_));
 sky130_fd_sc_hd__a21boi_2 _4498_ (.A1(_0615_),
    .A2(_0613_),
    .B1_N(_2688_),
    .Y(_0616_));
 sky130_fd_sc_hd__o21ai_2 _4499_ (.A1(_0616_),
    .A2(_2687_),
    .B1(_2685_),
    .Y(_0617_));
 sky130_fd_sc_hd__a21boi_2 _4500_ (.A1(_0612_),
    .A2(_0617_),
    .B1_N(_2682_),
    .Y(_0618_));
 sky130_fd_sc_hd__o21ai_2 _4501_ (.A1(_0618_),
    .A2(_2681_),
    .B1(_2679_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _4502_ (.A(_2673_),
    .B(_2676_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21oi_2 _4503_ (.A1(_0611_),
    .A2(_0619_),
    .B1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21o_1 _4504_ (.A1(_2673_),
    .A2(_2675_),
    .B1(_2672_),
    .X(_0622_));
 sky130_fd_sc_hd__o21ai_1 _4505_ (.A1(_0622_),
    .A2(_0621_),
    .B1(_2670_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2b_1 _4506_ (.A_N(_2669_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21o_1 _4507_ (.A1(_0624_),
    .A2(_2667_),
    .B1(_2666_),
    .X(_0625_));
 sky130_fd_sc_hd__a21o_1 _4508_ (.A1(_0625_),
    .A2(_2663_),
    .B1(_2662_),
    .X(_0626_));
 sky130_fd_sc_hd__and2_0 _4509_ (.A(_2654_),
    .B(_2657_),
    .X(_0627_));
 sky130_fd_sc_hd__a22o_1 _4510_ (.A1(_2654_),
    .A2(_2656_),
    .B1(_2659_),
    .B2(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__a311o_4 _4511_ (.A1(_2660_),
    .A2(_0627_),
    .A3(_0626_),
    .B1(_0628_),
    .C1(_2653_),
    .X(_0629_));
 sky130_fd_sc_hd__clkinv_4 _4512_ (.A(_0629_),
    .Y(_2868_));
 sky130_fd_sc_hd__o21ai_1 _4513_ (.A1(_2421_),
    .A2(_0321_),
    .B1(_2418_),
    .Y(_0630_));
 sky130_fd_sc_hd__a21oi_1 _4514_ (.A1(_0630_),
    .A2(_0326_),
    .B1(_0435_),
    .Y(_0631_));
 sky130_fd_sc_hd__o21a_1 _4515_ (.A1(_2405_),
    .A2(_0631_),
    .B1(_2540_),
    .X(_0632_));
 sky130_fd_sc_hd__nor3_1 _4516_ (.A(_2540_),
    .B(_2405_),
    .C(_0631_),
    .Y(_0633_));
 sky130_fd_sc_hd__nor2_2 _4517_ (.A(_0632_),
    .B(_0633_),
    .Y(_2618_));
 sky130_fd_sc_hd__inv_1 _4518_ (.A(_2487_),
    .Y(_0634_));
 sky130_fd_sc_hd__a21o_1 _4519_ (.A1(_2127_),
    .A2(_2497_),
    .B1(_2496_),
    .X(_0635_));
 sky130_fd_sc_hd__a21oi_1 _4520_ (.A1(_2491_),
    .A2(_0635_),
    .B1(_2490_),
    .Y(_0636_));
 sky130_fd_sc_hd__o21bai_1 _4521_ (.A1(_0634_),
    .A2(_0636_),
    .B1_N(_2486_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_2 _4522_ (.A1(_2484_),
    .A2(_0637_),
    .B1(_2483_),
    .Y(_0638_));
 sky130_fd_sc_hd__xnor2_2 _4523_ (.A(_2698_),
    .B(_0638_),
    .Y(_2699_));
 sky130_fd_sc_hd__inv_1 _4524_ (.A(_2699_),
    .Y(_2841_));
 sky130_fd_sc_hd__inv_1 _4525_ (.A(_2636_),
    .Y(_0639_));
 sky130_fd_sc_hd__o21ai_0 _4526_ (.A1(_0639_),
    .A2(_0610_),
    .B1(_0591_),
    .Y(_0640_));
 sky130_fd_sc_hd__a21oi_2 _4527_ (.A1(_2632_),
    .A2(_0640_),
    .B1(_2631_),
    .Y(_0641_));
 sky130_fd_sc_hd__xnor2_2 _4528_ (.A(_2628_),
    .B(_0641_),
    .Y(_2822_));
 sky130_fd_sc_hd__xor2_4 _4529_ (.A(_2624_),
    .B(_0604_),
    .X(_2818_));
 sky130_fd_sc_hd__inv_1 _4530_ (.A(_2709_),
    .Y(_0642_));
 sky130_fd_sc_hd__a21o_1 _4531_ (.A1(_2136_),
    .A2(_2719_),
    .B1(_2718_),
    .X(_0643_));
 sky130_fd_sc_hd__a21oi_1 _4532_ (.A1(_2713_),
    .A2(_0643_),
    .B1(_2712_),
    .Y(_0644_));
 sky130_fd_sc_hd__o21bai_1 _4533_ (.A1(_0642_),
    .A2(_0644_),
    .B1_N(_2708_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21oi_2 _4534_ (.A1(_2705_),
    .A2(_0645_),
    .B1(_2704_),
    .Y(_0646_));
 sky130_fd_sc_hd__xnor2_2 _4535_ (.A(_2702_),
    .B(_0646_),
    .Y(_2721_));
 sky130_fd_sc_hd__inv_1 _4536_ (.A(_2721_),
    .Y(_3024_));
 sky130_fd_sc_hd__a2111oi_1 _4537_ (.A1(_2386_),
    .A2(_2389_),
    .B1(_2531_),
    .C1(_2381_),
    .D1(_2385_),
    .Y(_0647_));
 sky130_fd_sc_hd__nor3_1 _4538_ (.A(_2382_),
    .B(_2381_),
    .C(_2531_),
    .Y(_0648_));
 sky130_fd_sc_hd__o31ai_1 _4539_ (.A1(_0533_),
    .A2(_0647_),
    .A3(_0648_),
    .B1(_0535_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _4540_ (.A1(_2580_),
    .A2(_0649_),
    .B1(_2579_),
    .X(_0650_));
 sky130_fd_sc_hd__nor2_1 _4541_ (.A(_0421_),
    .B(_0533_),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_2580_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nor2_1 _4543_ (.A(_0272_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_1 _4544_ (.A(_0650_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__xnor2_2 _4545_ (.A(_2726_),
    .B(_0654_),
    .Y(_2744_));
 sky130_fd_sc_hd__nor2b_1 _4546_ (.A(_2586_),
    .B_N(_0426_),
    .Y(_0655_));
 sky130_fd_sc_hd__a31oi_1 _4547_ (.A1(_0293_),
    .A2(_0537_),
    .A3(_0655_),
    .B1(_0159_),
    .Y(_0656_));
 sky130_fd_sc_hd__xnor2_1 _4548_ (.A(_2744_),
    .B(_0656_),
    .Y(_2727_));
 sky130_fd_sc_hd__nor2b_1 _4549_ (.A(_0306_),
    .B_N(_0655_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _4550_ (.A(net2),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__xnor2_1 _4551_ (.A(_2581_),
    .B(_0658_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_2536_),
    .B(_2734_),
    .Y(_0659_));
 sky130_fd_sc_hd__a21oi_1 _4553_ (.A1(_2734_),
    .A2(_2535_),
    .B1(_2733_),
    .Y(_0660_));
 sky130_fd_sc_hd__o21ai_2 _4554_ (.A1(_0437_),
    .A2(_0659_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__xor2_4 _4555_ (.A(_2730_),
    .B(_0661_),
    .X(_2748_));
 sky130_fd_sc_hd__a21oi_1 _4556_ (.A1(_2726_),
    .A2(_0650_),
    .B1(_2725_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand4_1 _4557_ (.A(_2580_),
    .B(_2726_),
    .C(_0280_),
    .D(_0651_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_0662_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__xor2_4 _4559_ (.A(_2738_),
    .B(_0664_),
    .X(_2739_));
 sky130_fd_sc_hd__o21a_1 _4560_ (.A1(_2583_),
    .A2(_0551_),
    .B1(_2746_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_1 _4561_ (.A(_2745_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__xnor2_4 _4562_ (.A(_2742_),
    .B(_0666_),
    .Y(_2768_));
 sky130_fd_sc_hd__a21boi_0 _4563_ (.A1(_2592_),
    .A2(_0562_),
    .B1_N(_0549_),
    .Y(_0667_));
 sky130_fd_sc_hd__o21bai_2 _4564_ (.A1(_0550_),
    .A2(_0667_),
    .B1_N(_2583_),
    .Y(_0668_));
 sky130_fd_sc_hd__xor2_4 _4565_ (.A(_2746_),
    .B(_0668_),
    .X(_2798_));
 sky130_fd_sc_hd__or4_1 _4566_ (.A(_2772_),
    .B(_0568_),
    .C(_0577_),
    .D(_2798_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(_0578_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__xor2_1 _4568_ (.A(_2768_),
    .B(_0670_),
    .X(_2747_));
 sky130_fd_sc_hd__o21ai_2 _4569_ (.A1(_2539_),
    .A2(_0632_),
    .B1(_2536_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2b_1 _4570_ (.A_N(_2535_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__xor2_2 _4571_ (.A(_2734_),
    .B(_0672_),
    .X(_2752_));
 sky130_fd_sc_hd__or3_1 _4572_ (.A(_0580_),
    .B(_2772_),
    .C(_0577_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(_0578_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__xor2_1 _4574_ (.A(_2798_),
    .B(_0674_),
    .X(_2751_));
 sky130_fd_sc_hd__o21ai_1 _4575_ (.A1(_2615_),
    .A2(_0603_),
    .B1(_2754_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(_2750_),
    .B(_2753_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _4577_ (.A(_2615_),
    .B(_2753_),
    .Y(_0677_));
 sky130_fd_sc_hd__o21ai_1 _4578_ (.A1(_2754_),
    .A2(_2753_),
    .B1(_2750_),
    .Y(_0678_));
 sky130_fd_sc_hd__a31oi_2 _4579_ (.A1(_0600_),
    .A2(_0602_),
    .A3(_0677_),
    .B1(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__a21oi_4 _4580_ (.A1(_0675_),
    .A2(_0676_),
    .B1(_0679_),
    .Y(_2806_));
 sky130_fd_sc_hd__and4_1 _4581_ (.A(_0012_),
    .B(_0053_),
    .C(_0171_),
    .D(_0214_),
    .X(_0680_));
 sky130_fd_sc_hd__nor4_2 _4582_ (.A(_0012_),
    .B(_0064_),
    .C(_0078_),
    .D(_0177_),
    .Y(_0681_));
 sky130_fd_sc_hd__o22ai_4 _4583_ (.A1(_0257_),
    .A2(_0258_),
    .B1(_0680_),
    .B2(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o211ai_2 _4584_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0251_),
    .C1(_0252_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor4_2 _4585_ (.A(_2566_),
    .B(_2574_),
    .C(_0682_),
    .D(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__xnor2_1 _4586_ (.A(_0032_),
    .B(_2087_),
    .Y(_0685_));
 sky130_fd_sc_hd__nor4_1 _4587_ (.A(_2088_),
    .B(_0025_),
    .C(_0113_),
    .D(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_1 _4588_ (.A(_0013_),
    .B(_0105_),
    .Y(_0687_));
 sky130_fd_sc_hd__a21oi_4 _4589_ (.A1(_0013_),
    .A2(_0686_),
    .B1(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nor4_2 _4590_ (.A(net16),
    .B(_2558_),
    .C(_2562_),
    .D(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__nor2_1 _4591_ (.A(_0226_),
    .B(_0439_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand4_1 _4592_ (.A(_0245_),
    .B(_0246_),
    .C(_0448_),
    .D(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_0229_),
    .B(_0448_),
    .Y(_0692_));
 sky130_fd_sc_hd__a31oi_1 _4594_ (.A1(_0451_),
    .A2(_0452_),
    .A3(_0692_),
    .B1(_0439_),
    .Y(_0693_));
 sky130_fd_sc_hd__nor3_1 _4595_ (.A(_2547_),
    .B(_0012_),
    .C(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__nor2_1 _4596_ (.A(_0450_),
    .B(_0491_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor3_1 _4597_ (.A(_2550_),
    .B(_2542_),
    .C(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _4598_ (.A(_2510_),
    .B(_2550_),
    .Y(_0697_));
 sky130_fd_sc_hd__o21ai_0 _4599_ (.A1(_2551_),
    .A2(_2550_),
    .B1(_0439_),
    .Y(_0698_));
 sky130_fd_sc_hd__a21oi_1 _4600_ (.A1(_0492_),
    .A2(_0697_),
    .B1(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_2542_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__a31oi_1 _4602_ (.A1(_0404_),
    .A2(_0407_),
    .A3(_0696_),
    .B1(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a22oi_2 _4603_ (.A1(_0691_),
    .A2(_0694_),
    .B1(_0701_),
    .B2(_0012_),
    .Y(_0702_));
 sky130_fd_sc_hd__xnor2_2 _4604_ (.A(_0478_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _4605_ (.A(net4),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__and2_0 _4606_ (.A(net4),
    .B(_0703_),
    .X(_0705_));
 sky130_fd_sc_hd__nand3_1 _4607_ (.A(_2580_),
    .B(_2726_),
    .C(_0651_),
    .Y(_0706_));
 sky130_fd_sc_hd__o21ai_0 _4608_ (.A1(_0272_),
    .A2(_0706_),
    .B1(_0662_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_1 _4609_ (.A1(_2738_),
    .A2(_0707_),
    .B1(_2737_),
    .Y(_0708_));
 sky130_fd_sc_hd__xnor3_1 _4610_ (.A(_0478_),
    .B(_0486_),
    .C(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__a2111oi_4 _4611_ (.A1(_0684_),
    .A2(_0689_),
    .B1(_0704_),
    .C1(_0705_),
    .D1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__and3_1 _4612_ (.A(_0709_),
    .B(_0684_),
    .C(_0689_),
    .X(_0711_));
 sky130_fd_sc_hd__o21a_1 _4613_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0709_),
    .X(_0712_));
 sky130_fd_sc_hd__or3_4 _4614_ (.A(_0710_),
    .B(_0711_),
    .C(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__inv_1 _4615_ (.A(_2744_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_1 _4616_ (.A(_0537_),
    .B(_0714_),
    .C(_0657_),
    .Y(_0715_));
 sky130_fd_sc_hd__buf_8 _4617_ (.A(_0295_),
    .X(_2124_));
 sky130_fd_sc_hd__o21ai_0 _4618_ (.A1(_2739_),
    .A2(_0715_),
    .B1(net23),
    .Y(_0716_));
 sky130_fd_sc_hd__o31ai_2 _4619_ (.A1(_0710_),
    .A2(_0711_),
    .A3(_0712_),
    .B1(net3),
    .Y(_0717_));
 sky130_fd_sc_hd__o21a_1 _4620_ (.A1(_0713_),
    .A2(_0716_),
    .B1(_0717_),
    .X(_2755_));
 sky130_fd_sc_hd__nor3_1 _4621_ (.A(_0710_),
    .B(_0711_),
    .C(_0712_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor2_1 _4622_ (.A(_2744_),
    .B(_2739_),
    .Y(_0719_));
 sky130_fd_sc_hd__a41o_1 _4623_ (.A1(_0293_),
    .A2(_0537_),
    .A3(_0655_),
    .A4(_0719_),
    .B1(net3),
    .X(_0720_));
 sky130_fd_sc_hd__xnor2_1 _4624_ (.A(_0718_),
    .B(_0720_),
    .Y(_2763_));
 sky130_fd_sc_hd__a31oi_1 _4625_ (.A1(_0537_),
    .A2(_0714_),
    .A3(_0657_),
    .B1(_0159_),
    .Y(_0721_));
 sky130_fd_sc_hd__xnor2_1 _4626_ (.A(_2739_),
    .B(_0721_),
    .Y(_2759_));
 sky130_fd_sc_hd__nor3_1 _4627_ (.A(_2535_),
    .B(_2729_),
    .C(_2733_),
    .Y(_0722_));
 sky130_fd_sc_hd__nor3_1 _4628_ (.A(_2734_),
    .B(_2729_),
    .C(_2733_),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _4629_ (.A(_2730_),
    .B(_2729_),
    .Y(_0724_));
 sky130_fd_sc_hd__a211oi_4 _4630_ (.A1(_0671_),
    .A2(_0722_),
    .B1(_0723_),
    .C1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21o_1 _4631_ (.A1(_2762_),
    .A2(_0725_),
    .B1(_2761_),
    .X(_0726_));
 sky130_fd_sc_hd__a21oi_2 _4632_ (.A1(_2766_),
    .A2(_0726_),
    .B1(_2765_),
    .Y(_0727_));
 sky130_fd_sc_hd__xnor2_4 _4633_ (.A(_2758_),
    .B(_0727_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21o_1 _4634_ (.A1(_2730_),
    .A2(_0661_),
    .B1(_2729_),
    .X(_0728_));
 sky130_fd_sc_hd__a21oi_4 _4635_ (.A1(_2762_),
    .A2(_0728_),
    .B1(_2761_),
    .Y(_0729_));
 sky130_fd_sc_hd__xnor2_4 _4636_ (.A(_2766_),
    .B(_0729_),
    .Y(_2928_));
 sky130_fd_sc_hd__inv_1 _4637_ (.A(_2762_),
    .Y(_0730_));
 sky130_fd_sc_hd__xnor2_4 _4638_ (.A(_0730_),
    .B(_0725_),
    .Y(_2932_));
 sky130_fd_sc_hd__inv_1 _4639_ (.A(_2788_),
    .Y(_0731_));
 sky130_fd_sc_hd__inv_1 _4640_ (.A(_2796_),
    .Y(_0732_));
 sky130_fd_sc_hd__inv_1 _4641_ (.A(_2484_),
    .Y(_0733_));
 sky130_fd_sc_hd__o21bai_1 _4642_ (.A1(_0733_),
    .A2(_0353_),
    .B1_N(_2483_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_2 _4643_ (.A1(_2698_),
    .A2(_0734_),
    .B1(_2697_),
    .Y(_0735_));
 sky130_fd_sc_hd__o21bai_1 _4644_ (.A1(_0732_),
    .A2(_0735_),
    .B1_N(_2795_),
    .Y(_0736_));
 sky130_fd_sc_hd__a21oi_1 _4645_ (.A1(_2792_),
    .A2(_0736_),
    .B1(_2791_),
    .Y(_0737_));
 sky130_fd_sc_hd__o21bai_1 _4646_ (.A1(_0731_),
    .A2(_0737_),
    .B1_N(_2787_),
    .Y(_0738_));
 sky130_fd_sc_hd__a21oi_2 _4647_ (.A1(_2784_),
    .A2(_0738_),
    .B1(_2783_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(_2804_),
    .B(_2780_),
    .Y(_0740_));
 sky130_fd_sc_hd__a21oi_1 _4649_ (.A1(_2804_),
    .A2(_2779_),
    .B1(_2803_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21ai_2 _4650_ (.A1(_0739_),
    .A2(_0740_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__a21o_1 _4651_ (.A1(_2776_),
    .A2(_0742_),
    .B1(_2773_),
    .X(_0743_));
 sky130_fd_sc_hd__a21oi_1 _4652_ (.A1(_2800_),
    .A2(_0743_),
    .B1(_2799_),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_2 _4653_ (.A(_2770_),
    .B(_0744_),
    .Y(_2948_));
 sky130_fd_sc_hd__nand2_1 _4654_ (.A(_2804_),
    .B(_2776_),
    .Y(_0745_));
 sky130_fd_sc_hd__inv_1 _4655_ (.A(_2698_),
    .Y(_0746_));
 sky130_fd_sc_hd__o21bai_1 _4656_ (.A1(_0746_),
    .A2(_0638_),
    .B1_N(_2697_),
    .Y(_0747_));
 sky130_fd_sc_hd__a211oi_1 _4657_ (.A1(_2796_),
    .A2(_0747_),
    .B1(_2795_),
    .C1(_2791_),
    .Y(_0748_));
 sky130_fd_sc_hd__o21ai_0 _4658_ (.A1(_2792_),
    .A2(_2791_),
    .B1(_2788_),
    .Y(_0749_));
 sky130_fd_sc_hd__o21bai_2 _4659_ (.A1(_0748_),
    .A2(_0749_),
    .B1_N(_2787_),
    .Y(_0750_));
 sky130_fd_sc_hd__a21o_1 _4660_ (.A1(_2784_),
    .A2(_0750_),
    .B1(_2783_),
    .X(_0751_));
 sky130_fd_sc_hd__a21oi_2 _4661_ (.A1(_2780_),
    .A2(_0751_),
    .B1(_2779_),
    .Y(_0752_));
 sky130_fd_sc_hd__a21oi_1 _4662_ (.A1(_2774_),
    .A2(_2803_),
    .B1(_2773_),
    .Y(_0753_));
 sky130_fd_sc_hd__o21ai_1 _4663_ (.A1(_0745_),
    .A2(_0752_),
    .B1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__xor2_2 _4664_ (.A(_2800_),
    .B(_0754_),
    .X(_2974_));
 sky130_fd_sc_hd__xor2_4 _4665_ (.A(_2776_),
    .B(_0742_),
    .X(_2952_));
 sky130_fd_sc_hd__xnor2_2 _4666_ (.A(_2804_),
    .B(_0752_),
    .Y(_2978_));
 sky130_fd_sc_hd__xnor2_2 _4667_ (.A(_2780_),
    .B(_0739_),
    .Y(_2958_));
 sky130_fd_sc_hd__xor2_2 _4668_ (.A(_2784_),
    .B(_0750_),
    .X(_2962_));
 sky130_fd_sc_hd__a21oi_1 _4669_ (.A1(_2796_),
    .A2(_0747_),
    .B1(_2795_),
    .Y(_0755_));
 sky130_fd_sc_hd__xnor2_2 _4670_ (.A(_2792_),
    .B(_0755_),
    .Y(_2970_));
 sky130_fd_sc_hd__xnor2_2 _4671_ (.A(_2788_),
    .B(_0737_),
    .Y(_2966_));
 sky130_fd_sc_hd__or2_0 _4672_ (.A(_2970_),
    .B(_2966_),
    .X(_0756_));
 sky130_fd_sc_hd__or2_0 _4673_ (.A(_2962_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__xnor2_2 _4674_ (.A(_2796_),
    .B(_0735_),
    .Y(_2896_));
 sky130_fd_sc_hd__or3_1 _4675_ (.A(_2499_),
    .B(_2699_),
    .C(_2896_),
    .X(_0758_));
 sky130_fd_sc_hd__or3_1 _4676_ (.A(_2958_),
    .B(_0757_),
    .C(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__or3_1 _4677_ (.A(_2952_),
    .B(_2978_),
    .C(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__o31a_1 _4678_ (.A1(_2948_),
    .A2(_2974_),
    .A3(_0760_),
    .B1(net13),
    .X(_0761_));
 sky130_fd_sc_hd__nand2b_1 _4679_ (.A_N(_2417_),
    .B(_0630_),
    .Y(_0762_));
 sky130_fd_sc_hd__a21oi_2 _4680_ (.A1(_2414_),
    .A2(_0762_),
    .B1(_2413_),
    .Y(_0763_));
 sky130_fd_sc_hd__xnor2_4 _4681_ (.A(_2410_),
    .B(_0763_),
    .Y(_2626_));
 sky130_fd_sc_hd__or3_1 _4682_ (.A(_2630_),
    .B(_2634_),
    .C(_2638_),
    .X(_0764_));
 sky130_fd_sc_hd__nor4_1 _4683_ (.A(_2622_),
    .B(_2618_),
    .C(_2626_),
    .D(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_0438_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__or3_1 _4685_ (.A(_2748_),
    .B(_2752_),
    .C(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__nor4_1 _4686_ (.A(_2944_),
    .B(_2928_),
    .C(_2932_),
    .D(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_2758_),
    .B(_2766_),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_1 _4688_ (.A1(_2758_),
    .A2(_2765_),
    .B1(_2757_),
    .Y(_0770_));
 sky130_fd_sc_hd__o21ai_2 _4689_ (.A1(_0729_),
    .A2(_0769_),
    .B1(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__o211ai_4 _4690_ (.A1(_0713_),
    .A2(_0720_),
    .B1(_0771_),
    .C1(_0717_),
    .Y(_0772_));
 sky130_fd_sc_hd__nor4b_1 _4691_ (.A(_0710_),
    .B(_0711_),
    .C(_0712_),
    .D_N(_0720_),
    .Y(_0773_));
 sky130_fd_sc_hd__a211o_2 _4692_ (.A1(net18),
    .A2(_0713_),
    .B1(_0773_),
    .C1(_0771_),
    .X(_0774_));
 sky130_fd_sc_hd__a21o_1 _4693_ (.A1(_2564_),
    .A2(_0527_),
    .B1(_2563_),
    .X(_0775_));
 sky130_fd_sc_hd__a21oi_2 _4694_ (.A1(_2560_),
    .A2(_0775_),
    .B1(_2559_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor3_1 _4695_ (.A(net16),
    .B(_2736_),
    .C(_2724_),
    .Y(_0777_));
 sky130_fd_sc_hd__xnor2_1 _4696_ (.A(net16),
    .B(_0478_),
    .Y(_0778_));
 sky130_fd_sc_hd__xnor2_1 _4697_ (.A(_0486_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__a31oi_2 _4698_ (.A1(_0496_),
    .A2(_0500_),
    .A3(_0777_),
    .B1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__xnor2_2 _4699_ (.A(_0703_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__xor2_4 _4700_ (.A(_0776_),
    .B(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__a21oi_2 _4701_ (.A1(_0772_),
    .A2(_0774_),
    .B1(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__and3_1 _4702_ (.A(_0772_),
    .B(_0774_),
    .C(_0782_),
    .X(_0784_));
 sky130_fd_sc_hd__or4_2 _4703_ (.A(_2665_),
    .B(_0768_),
    .C(_0783_),
    .D(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__o21ai_2 _4704_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_2665_),
    .Y(_0786_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_2769_),
    .B(_2799_),
    .Y(_0787_));
 sky130_fd_sc_hd__o211ai_1 _4706_ (.A1(_0745_),
    .A2(_0752_),
    .B1(_0753_),
    .C1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__or3_1 _4707_ (.A(_2800_),
    .B(_2769_),
    .C(_2799_),
    .X(_0789_));
 sky130_fd_sc_hd__o211ai_1 _4708_ (.A1(_2770_),
    .A2(_2769_),
    .B1(_0788_),
    .C1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor4_1 _4709_ (.A(_2764_),
    .B(_2760_),
    .C(_2728_),
    .D(_2732_),
    .Y(_0791_));
 sky130_fd_sc_hd__xnor2_2 _4710_ (.A(_2270_),
    .B(_0299_),
    .Y(_2416_));
 sky130_fd_sc_hd__or3_1 _4711_ (.A(_2420_),
    .B(_2424_),
    .C(_2416_),
    .X(_0792_));
 sky130_fd_sc_hd__or3_1 _4712_ (.A(_2412_),
    .B(_2408_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__or4_1 _4713_ (.A(_2404_),
    .B(_2534_),
    .C(_2538_),
    .D(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_1 _4714_ (.A(_2756_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__a21oi_2 _4715_ (.A1(_0791_),
    .A2(_0795_),
    .B1(net3),
    .Y(_0796_));
 sky130_fd_sc_hd__mux2i_4 _4716_ (.A0(net3),
    .A1(_0796_),
    .S(_0782_),
    .Y(_0797_));
 sky130_fd_sc_hd__a21o_1 _4717_ (.A1(_2746_),
    .A2(_0668_),
    .B1(_2745_),
    .X(_0798_));
 sky130_fd_sc_hd__a21oi_2 _4718_ (.A1(_2742_),
    .A2(_0798_),
    .B1(_2741_),
    .Y(_0799_));
 sky130_fd_sc_hd__xnor2_4 _4719_ (.A(_0713_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor3_1 _4720_ (.A(_0790_),
    .B(_0797_),
    .C(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__a21oi_4 _4721_ (.A1(_0785_),
    .A2(_0786_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__and3_2 _4722_ (.A(_0785_),
    .B(_0786_),
    .C(_0801_),
    .X(_0803_));
 sky130_fd_sc_hd__or2_0 _4723_ (.A(_0802_),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__xor2_1 _4724_ (.A(_0761_),
    .B(_0804_),
    .X(_2805_));
 sky130_fd_sc_hd__inv_1 _4725_ (.A(_2628_),
    .Y(_0805_));
 sky130_fd_sc_hd__o21ai_0 _4726_ (.A1(_0805_),
    .A2(_0641_),
    .B1(_0590_),
    .Y(_0806_));
 sky130_fd_sc_hd__a21oi_1 _4727_ (.A1(_2624_),
    .A2(_0806_),
    .B1(_2623_),
    .Y(_0807_));
 sky130_fd_sc_hd__nor2b_1 _4728_ (.A(_0807_),
    .B_N(_2620_),
    .Y(_0808_));
 sky130_fd_sc_hd__o21a_1 _4729_ (.A1(_2619_),
    .A2(_0808_),
    .B1(_2616_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_2 _4730_ (.A(_2615_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__xnor2_4 _4731_ (.A(_2754_),
    .B(_0810_),
    .Y(_2810_));
 sky130_fd_sc_hd__buf_6 _4732_ (.A(_0629_),
    .X(_2852_));
 sky130_fd_sc_hd__nand2b_1 _4733_ (.A_N(_2896_),
    .B(_2843_),
    .Y(_0811_));
 sky130_fd_sc_hd__nor4_1 _4734_ (.A(_2978_),
    .B(_2958_),
    .C(_0757_),
    .D(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nor2_1 _4735_ (.A(_2974_),
    .B(_2952_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand2_1 _4736_ (.A(_0812_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(net12),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__xor2_1 _4738_ (.A(_2948_),
    .B(_0815_),
    .X(_2809_));
 sky130_fd_sc_hd__buf_2 _4739_ (.A(_0629_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_0816_),
    .B(_0760_),
    .Y(_0817_));
 sky130_fd_sc_hd__xor2_1 _4741_ (.A(_2974_),
    .B(_0817_),
    .X(_2847_));
 sky130_fd_sc_hd__nor2_1 _4742_ (.A(net1),
    .B(_0812_),
    .Y(_0818_));
 sky130_fd_sc_hd__xnor2_1 _4743_ (.A(_2952_),
    .B(_0818_),
    .Y(_2813_));
 sky130_fd_sc_hd__nand2_1 _4744_ (.A(_0816_),
    .B(_0759_),
    .Y(_0819_));
 sky130_fd_sc_hd__xor2_1 _4745_ (.A(_2978_),
    .B(_0819_),
    .X(_2817_));
 sky130_fd_sc_hd__o21ai_0 _4746_ (.A1(_0757_),
    .A2(_0811_),
    .B1(_0816_),
    .Y(_0820_));
 sky130_fd_sc_hd__xor2_1 _4747_ (.A(_2958_),
    .B(_0820_),
    .X(_2821_));
 sky130_fd_sc_hd__o21ai_0 _4748_ (.A1(_0756_),
    .A2(_0758_),
    .B1(_0816_),
    .Y(_0821_));
 sky130_fd_sc_hd__xor2_1 _4749_ (.A(_2962_),
    .B(_0821_),
    .X(_2825_));
 sky130_fd_sc_hd__o21ai_0 _4750_ (.A1(_2970_),
    .A2(_0811_),
    .B1(_0816_),
    .Y(_0822_));
 sky130_fd_sc_hd__xor2_1 _4751_ (.A(_2966_),
    .B(_0822_),
    .X(_2829_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_0816_),
    .B(_0758_),
    .Y(_0823_));
 sky130_fd_sc_hd__xor2_1 _4753_ (.A(_2970_),
    .B(_0823_),
    .X(_2833_));
 sky130_fd_sc_hd__nor2_1 _4754_ (.A(_2843_),
    .B(_2868_),
    .Y(_0824_));
 sky130_fd_sc_hd__xnor2_1 _4755_ (.A(_2896_),
    .B(_0824_),
    .Y(_2837_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_2844_),
    .B(_0816_),
    .Y(_0825_));
 sky130_fd_sc_hd__o21ai_1 _4757_ (.A1(_0816_),
    .A2(_2841_),
    .B1(_0825_),
    .Y(_2141_));
 sky130_fd_sc_hd__inv_1 _4758_ (.A(_2141_),
    .Y(_2145_));
 sky130_fd_sc_hd__inv_1 _4759_ (.A(_2823_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_1 _4760_ (.A(_2831_),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_1 _4761_ (.A(_2839_),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2b_1 _4762_ (.A(_2140_),
    .B_N(_2846_),
    .Y(_0829_));
 sky130_fd_sc_hd__o21ai_1 _4763_ (.A1(_2845_),
    .A2(_0829_),
    .B1(_2840_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21boi_0 _4764_ (.A1(_0828_),
    .A2(_0830_),
    .B1_N(_2836_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21ai_1 _4765_ (.A1(_2835_),
    .A2(_0831_),
    .B1(_2832_),
    .Y(_0832_));
 sky130_fd_sc_hd__a21boi_1 _4766_ (.A1(_0827_),
    .A2(_0832_),
    .B1_N(_2828_),
    .Y(_0833_));
 sky130_fd_sc_hd__o21ai_1 _4767_ (.A1(_2827_),
    .A2(_0833_),
    .B1(_2824_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21boi_1 _4768_ (.A1(_0826_),
    .A2(_0834_),
    .B1_N(_2820_),
    .Y(_0835_));
 sky130_fd_sc_hd__o21ai_0 _4769_ (.A1(_2819_),
    .A2(_0835_),
    .B1(_2816_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2b_1 _4770_ (.A_N(_2815_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a21o_1 _4771_ (.A1(_2850_),
    .A2(_0837_),
    .B1(_2849_),
    .X(_0838_));
 sky130_fd_sc_hd__a21o_2 _4772_ (.A1(_2812_),
    .A2(_0838_),
    .B1(_2811_),
    .X(_0839_));
 sky130_fd_sc_hd__xor2_4 _4773_ (.A(_2808_),
    .B(_0839_),
    .X(_3034_));
 sky130_fd_sc_hd__xor2_2 _4774_ (.A(_2850_),
    .B(_0837_),
    .X(_2992_));
 sky130_fd_sc_hd__nand2_1 _4775_ (.A(_0826_),
    .B(_0834_),
    .Y(_0840_));
 sky130_fd_sc_hd__nor2_1 _4776_ (.A(_2820_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nor2_2 _4777_ (.A(_0835_),
    .B(_0841_),
    .Y(_3000_));
 sky130_fd_sc_hd__inv_1 _4778_ (.A(_2827_),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_1 _4779_ (.A(_2835_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2b_1 _4780_ (.A(_2143_),
    .B_N(_2840_),
    .Y(_0844_));
 sky130_fd_sc_hd__o21ai_0 _4781_ (.A1(_2839_),
    .A2(_0844_),
    .B1(_2836_),
    .Y(_0845_));
 sky130_fd_sc_hd__a21boi_0 _4782_ (.A1(_0843_),
    .A2(_0845_),
    .B1_N(_2832_),
    .Y(_0846_));
 sky130_fd_sc_hd__o21ai_0 _4783_ (.A1(_2831_),
    .A2(_0846_),
    .B1(_2828_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21boi_0 _4784_ (.A1(_0842_),
    .A2(_0847_),
    .B1_N(_2824_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_0842_),
    .B(_0847_),
    .Y(_0849_));
 sky130_fd_sc_hd__nor2_1 _4786_ (.A(_2824_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_1 _4787_ (.A(_0848_),
    .B(_0850_),
    .Y(_3004_));
 sky130_fd_sc_hd__inv_1 _4788_ (.A(_3004_),
    .Y(_2919_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_0827_),
    .B(_0832_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_1 _4790_ (.A(_2828_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_2 _4791_ (.A(_0833_),
    .B(_0852_),
    .Y(_3008_));
 sky130_fd_sc_hd__inv_1 _4792_ (.A(_3008_),
    .Y(_2918_));
 sky130_fd_sc_hd__inv_1 _4793_ (.A(_2863_),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_1 _4794_ (.A(_2870_),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_1 _4795_ (.A(_2876_),
    .Y(_0855_));
 sky130_fd_sc_hd__inv_1 _4796_ (.A(_2882_),
    .Y(_0856_));
 sky130_fd_sc_hd__inv_1 _4797_ (.A(_2888_),
    .Y(_0857_));
 sky130_fd_sc_hd__a21o_1 _4798_ (.A1(_2894_),
    .A2(net62),
    .B1(_2893_),
    .X(_0858_));
 sky130_fd_sc_hd__a21oi_2 _4799_ (.A1(_0858_),
    .A2(_2891_),
    .B1(_2890_),
    .Y(_0859_));
 sky130_fd_sc_hd__inv_1 _4800_ (.A(_2887_),
    .Y(_0860_));
 sky130_fd_sc_hd__o21ai_1 _4801_ (.A1(_0857_),
    .A2(_0859_),
    .B1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__a21oi_2 _4802_ (.A1(_0861_),
    .A2(_2885_),
    .B1(_2884_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21bai_1 _4803_ (.A1(_0856_),
    .A2(_0862_),
    .B1_N(_2881_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_2 _4804_ (.A1(_0863_),
    .A2(_2879_),
    .B1(_2878_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21bai_1 _4805_ (.A1(_0864_),
    .A2(_0855_),
    .B1_N(_2875_),
    .Y(_0865_));
 sky130_fd_sc_hd__a21oi_2 _4806_ (.A1(_0865_),
    .A2(_2873_),
    .B1(_2872_),
    .Y(_0866_));
 sky130_fd_sc_hd__o21bai_1 _4807_ (.A1(_0854_),
    .A2(_0866_),
    .B1_N(_2869_),
    .Y(_0867_));
 sky130_fd_sc_hd__a21oi_2 _4808_ (.A1(_0867_),
    .A2(_2866_),
    .B1(_2865_),
    .Y(_0868_));
 sky130_fd_sc_hd__o21bai_1 _4809_ (.A1(_0868_),
    .A2(_0853_),
    .B1_N(_2862_),
    .Y(_0869_));
 sky130_fd_sc_hd__a21oi_2 _4810_ (.A1(_0869_),
    .A2(_2860_),
    .B1(_2859_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_2854_),
    .B(_2857_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21oi_1 _4812_ (.A1(_2854_),
    .A2(_2856_),
    .B1(_2853_),
    .Y(_0872_));
 sky130_fd_sc_hd__o21ai_4 _4813_ (.A1(_0871_),
    .A2(_0870_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__clkinv_4 _4814_ (.A(_0873_),
    .Y(_3057_));
 sky130_fd_sc_hd__xnor2_2 _4815_ (.A(_2620_),
    .B(_0807_),
    .Y(_2814_));
 sky130_fd_sc_hd__inv_1 _4816_ (.A(_2705_),
    .Y(_0874_));
 sky130_fd_sc_hd__a21oi_1 _4817_ (.A1(_2713_),
    .A2(_2138_),
    .B1(_2712_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_0642_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__nor2_1 _4819_ (.A(_2708_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__o21bai_1 _4820_ (.A1(_0874_),
    .A2(_0877_),
    .B1_N(_2704_),
    .Y(_0878_));
 sky130_fd_sc_hd__a21oi_1 _4821_ (.A1(_2702_),
    .A2(_0878_),
    .B1(_2701_),
    .Y(_0879_));
 sky130_fd_sc_hd__xnor2_2 _4822_ (.A(_2898_),
    .B(_0879_),
    .Y(_2899_));
 sky130_fd_sc_hd__inv_1 _4823_ (.A(_2899_),
    .Y(_3023_));
 sky130_fd_sc_hd__inv_1 _4824_ (.A(_2819_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ai_0 _4825_ (.A1(_2823_),
    .A2(_0848_),
    .B1(_2820_),
    .Y(_0881_));
 sky130_fd_sc_hd__a21boi_1 _4826_ (.A1(_0880_),
    .A2(_0881_),
    .B1_N(_2816_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2_1 _4827_ (.A(_0880_),
    .B(_0881_),
    .Y(_0883_));
 sky130_fd_sc_hd__nor2_1 _4828_ (.A(_2816_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_2 _4829_ (.A(_0882_),
    .B(_0884_),
    .Y(_2996_));
 sky130_fd_sc_hd__inv_1 _4830_ (.A(_2849_),
    .Y(_0885_));
 sky130_fd_sc_hd__o21ai_0 _4831_ (.A1(_2815_),
    .A2(_0882_),
    .B1(_2850_),
    .Y(_0886_));
 sky130_fd_sc_hd__a21boi_1 _4832_ (.A1(_0885_),
    .A2(_0886_),
    .B1_N(_2812_),
    .Y(_0887_));
 sky130_fd_sc_hd__nand2_1 _4833_ (.A(_0885_),
    .B(_0886_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_1 _4834_ (.A(_2812_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_2 _4835_ (.A(_0887_),
    .B(_0889_),
    .Y(_2986_));
 sky130_fd_sc_hd__inv_1 _4836_ (.A(_2909_),
    .Y(_0890_));
 sky130_fd_sc_hd__inv_1 _4837_ (.A(_2913_),
    .Y(_0891_));
 sky130_fd_sc_hd__a21oi_1 _4838_ (.A1(_2148_),
    .A2(_2917_),
    .B1(_2916_),
    .Y(_0892_));
 sky130_fd_sc_hd__nor2_1 _4839_ (.A(_0891_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_1 _4840_ (.A(_2912_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__o21bai_1 _4841_ (.A1(_0890_),
    .A2(_0894_),
    .B1_N(_2908_),
    .Y(_0895_));
 sky130_fd_sc_hd__a21oi_2 _4842_ (.A1(_2905_),
    .A2(_0895_),
    .B1(_2904_),
    .Y(_0896_));
 sky130_fd_sc_hd__xnor2_4 _4843_ (.A(_2902_),
    .B(_0896_),
    .Y(_2925_));
 sky130_fd_sc_hd__inv_1 _4844_ (.A(_2925_),
    .Y(_3192_));
 sky130_fd_sc_hd__o211a_1 _4845_ (.A1(_2768_),
    .A2(_0669_),
    .B1(_0800_),
    .C1(net6),
    .X(_0897_));
 sky130_fd_sc_hd__o21ai_0 _4846_ (.A1(_2768_),
    .A2(_0669_),
    .B1(net6),
    .Y(_0898_));
 sky130_fd_sc_hd__nor2_1 _4847_ (.A(_0800_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__mux2i_4 _4848_ (.A0(_0897_),
    .A1(_0899_),
    .S(_0797_),
    .Y(_0900_));
 sky130_fd_sc_hd__nor2_1 _4849_ (.A(net6),
    .B(_0800_),
    .Y(_0901_));
 sky130_fd_sc_hd__and2_0 _4850_ (.A(_2665_),
    .B(_0800_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2i_4 _4851_ (.A0(_0901_),
    .A1(_0902_),
    .S(_0797_),
    .Y(_0903_));
 sky130_fd_sc_hd__and2_0 _4852_ (.A(_0900_),
    .B(_0903_),
    .X(_2927_));
 sky130_fd_sc_hd__xnor2_1 _4853_ (.A(_0797_),
    .B(_0800_),
    .Y(_0904_));
 sky130_fd_sc_hd__o31ai_2 _4854_ (.A1(_2768_),
    .A2(_2798_),
    .A3(_0673_),
    .B1(_0578_),
    .Y(_0905_));
 sky130_fd_sc_hd__xor2_1 _4855_ (.A(_0904_),
    .B(_0905_),
    .X(_2931_));
 sky130_fd_sc_hd__o21ai_0 _4856_ (.A1(_2749_),
    .A2(_0679_),
    .B1(_2934_),
    .Y(_0906_));
 sky130_fd_sc_hd__nand2b_1 _4857_ (.A_N(_2933_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__xnor2_2 _4858_ (.A(_2930_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__inv_1 _4859_ (.A(_0908_),
    .Y(_2936_));
 sky130_fd_sc_hd__o21ai_2 _4860_ (.A1(_0802_),
    .A2(_0803_),
    .B1(_0761_),
    .Y(_0909_));
 sky130_fd_sc_hd__or3_2 _4861_ (.A(net13),
    .B(_0802_),
    .C(_0803_),
    .X(_0910_));
 sky130_fd_sc_hd__and2_0 _4862_ (.A(_0909_),
    .B(_0910_),
    .X(_2935_));
 sky130_fd_sc_hd__nor3_1 _4863_ (.A(_2754_),
    .B(_2749_),
    .C(_2753_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_2750_),
    .B(_2749_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_1 _4865_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__o41ai_4 _4866_ (.A1(_2615_),
    .A2(_2749_),
    .A3(_2753_),
    .A4(_0809_),
    .B1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__xnor2_2 _4867_ (.A(_2934_),
    .B(_0914_),
    .Y(_2940_));
 sky130_fd_sc_hd__o211ai_1 _4868_ (.A1(_2948_),
    .A2(_0814_),
    .B1(_0804_),
    .C1(_0816_),
    .Y(_0915_));
 sky130_fd_sc_hd__and2_0 _4869_ (.A(_0910_),
    .B(_0915_),
    .X(_2939_));
 sky130_fd_sc_hd__a21o_1 _4870_ (.A1(_2942_),
    .A2(_2807_),
    .B1(_2941_),
    .X(_0916_));
 sky130_fd_sc_hd__a31oi_4 _4871_ (.A1(_2808_),
    .A2(_2942_),
    .A3(_0839_),
    .B1(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__xnor2_4 _4872_ (.A(_2938_),
    .B(_0917_),
    .Y(_2981_));
 sky130_fd_sc_hd__o21a_1 _4873_ (.A1(_0904_),
    .A2(_0905_),
    .B1(_0903_),
    .X(_2943_));
 sky130_fd_sc_hd__inv_1 _4874_ (.A(_2934_),
    .Y(_0918_));
 sky130_fd_sc_hd__o21bai_1 _4875_ (.A1(_0918_),
    .A2(_0914_),
    .B1_N(_2933_),
    .Y(_0919_));
 sky130_fd_sc_hd__a21oi_1 _4876_ (.A1(_2930_),
    .A2(_0919_),
    .B1(_2929_),
    .Y(_0920_));
 sky130_fd_sc_hd__xor2_1 _4877_ (.A(_2946_),
    .B(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__inv_1 _4878_ (.A(_0921_),
    .Y(_3117_));
 sky130_fd_sc_hd__inv_1 _4879_ (.A(_2956_),
    .Y(_0922_));
 sky130_fd_sc_hd__inv_1 _4880_ (.A(_2960_),
    .Y(_0923_));
 sky130_fd_sc_hd__inv_1 _4881_ (.A(_2968_),
    .Y(_0924_));
 sky130_fd_sc_hd__inv_1 _4882_ (.A(_2898_),
    .Y(_0925_));
 sky130_fd_sc_hd__o21bai_1 _4883_ (.A1(_0925_),
    .A2(_0879_),
    .B1_N(_2897_),
    .Y(_0926_));
 sky130_fd_sc_hd__a21oi_1 _4884_ (.A1(_2972_),
    .A2(_0926_),
    .B1(_2971_),
    .Y(_0927_));
 sky130_fd_sc_hd__o21bai_1 _4885_ (.A1(_0924_),
    .A2(_0927_),
    .B1_N(_2967_),
    .Y(_0928_));
 sky130_fd_sc_hd__a21oi_1 _4886_ (.A1(_2964_),
    .A2(_0928_),
    .B1(_2963_),
    .Y(_0929_));
 sky130_fd_sc_hd__o21bai_1 _4887_ (.A1(_0923_),
    .A2(_0929_),
    .B1_N(_2959_),
    .Y(_0930_));
 sky130_fd_sc_hd__a21oi_2 _4888_ (.A1(_2980_),
    .A2(_0930_),
    .B1(_2979_),
    .Y(_0931_));
 sky130_fd_sc_hd__o21bai_1 _4889_ (.A1(_0922_),
    .A2(_0931_),
    .B1_N(_2953_),
    .Y(_0932_));
 sky130_fd_sc_hd__a21oi_2 _4890_ (.A1(_2976_),
    .A2(_0932_),
    .B1(_2975_),
    .Y(_0933_));
 sky130_fd_sc_hd__xnor2_4 _4891_ (.A(_2950_),
    .B(_0933_),
    .Y(_3126_));
 sky130_fd_sc_hd__inv_1 _4892_ (.A(_2964_),
    .Y(_0934_));
 sky130_fd_sc_hd__inv_1 _4893_ (.A(_2972_),
    .Y(_0935_));
 sky130_fd_sc_hd__inv_1 _4894_ (.A(_2702_),
    .Y(_0936_));
 sky130_fd_sc_hd__o21bai_1 _4895_ (.A1(_0936_),
    .A2(_0646_),
    .B1_N(_2701_),
    .Y(_0937_));
 sky130_fd_sc_hd__a21oi_2 _4896_ (.A1(_2898_),
    .A2(_0937_),
    .B1(_2897_),
    .Y(_0938_));
 sky130_fd_sc_hd__o21bai_1 _4897_ (.A1(_0935_),
    .A2(_0938_),
    .B1_N(_2971_),
    .Y(_0939_));
 sky130_fd_sc_hd__a21oi_1 _4898_ (.A1(_2968_),
    .A2(_0939_),
    .B1(_2967_),
    .Y(_0940_));
 sky130_fd_sc_hd__o21bai_1 _4899_ (.A1(_0934_),
    .A2(_0940_),
    .B1_N(_2963_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21oi_4 _4900_ (.A1(_2960_),
    .A2(_0941_),
    .B1(_2959_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(_2980_),
    .B(_2956_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21oi_2 _4902_ (.A1(_2954_),
    .A2(_2979_),
    .B1(_2953_),
    .Y(_0944_));
 sky130_fd_sc_hd__o21ai_4 _4903_ (.A1(_0942_),
    .A2(_0943_),
    .B1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__xor2_4 _4904_ (.A(_2976_),
    .B(_0945_),
    .X(_3130_));
 sky130_fd_sc_hd__xnor2_4 _4905_ (.A(_2956_),
    .B(_0931_),
    .Y(_3134_));
 sky130_fd_sc_hd__xnor2_4 _4906_ (.A(_2980_),
    .B(_0942_),
    .Y(_3152_));
 sky130_fd_sc_hd__xnor2_2 _4907_ (.A(_2960_),
    .B(_0929_),
    .Y(_3138_));
 sky130_fd_sc_hd__xnor2_2 _4908_ (.A(_2964_),
    .B(_0940_),
    .Y(_3142_));
 sky130_fd_sc_hd__xnor2_2 _4909_ (.A(_2968_),
    .B(_0927_),
    .Y(_3146_));
 sky130_fd_sc_hd__and2_0 _4910_ (.A(_0772_),
    .B(_0774_),
    .X(_0946_));
 sky130_fd_sc_hd__a21o_1 _4911_ (.A1(_2946_),
    .A2(_2929_),
    .B1(_2945_),
    .X(_0947_));
 sky130_fd_sc_hd__a31oi_1 _4912_ (.A1(_2930_),
    .A2(_2946_),
    .A3(_0907_),
    .B1(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__xor3_1 _4913_ (.A(_0946_),
    .B(_0782_),
    .C(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__a21oi_4 _4914_ (.A1(_0900_),
    .A2(_0903_),
    .B1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__and3_2 _4915_ (.A(_0900_),
    .B(_0903_),
    .C(_0949_),
    .X(_0951_));
 sky130_fd_sc_hd__or3_2 _4916_ (.A(net13),
    .B(_0950_),
    .C(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__or3_1 _4917_ (.A(_2826_),
    .B(_2830_),
    .C(_2822_),
    .X(_0953_));
 sky130_fd_sc_hd__or3_1 _4918_ (.A(_2818_),
    .B(_2814_),
    .C(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__or3_1 _4919_ (.A(_2848_),
    .B(_2810_),
    .C(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__nor3_1 _4920_ (.A(_2806_),
    .B(_2940_),
    .C(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__a31oi_2 _4921_ (.A1(_0908_),
    .A2(_0921_),
    .A3(_0956_),
    .B1(net1),
    .Y(_0957_));
 sky130_fd_sc_hd__o21ai_2 _4922_ (.A1(_0950_),
    .A2(_0951_),
    .B1(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand3_1 _4923_ (.A(_2950_),
    .B(_2976_),
    .C(_0945_),
    .Y(_0959_));
 sky130_fd_sc_hd__a21oi_1 _4924_ (.A1(_2950_),
    .A2(_2975_),
    .B1(_2949_),
    .Y(_0960_));
 sky130_fd_sc_hd__nand2_1 _4925_ (.A(_0959_),
    .B(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__o21ai_2 _4926_ (.A1(_0802_),
    .A2(_0803_),
    .B1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__or3_1 _4927_ (.A(_0802_),
    .B(_0803_),
    .C(_0961_),
    .X(_0963_));
 sky130_fd_sc_hd__a22oi_4 _4928_ (.A1(_0952_),
    .A2(_0958_),
    .B1(_0962_),
    .B2(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__and4_2 _4929_ (.A(_0952_),
    .B(_0958_),
    .C(_0962_),
    .D(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_3024_),
    .B(_3023_),
    .Y(_0966_));
 sky130_fd_sc_hd__xnor2_4 _4931_ (.A(_2972_),
    .B(_0938_),
    .Y(_3082_));
 sky130_fd_sc_hd__nor2_1 _4932_ (.A(_3146_),
    .B(_3082_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand2b_1 _4933_ (.A_N(_3142_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__nor2_1 _4934_ (.A(_3138_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2b_1 _4935_ (.A_N(_3152_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__or4_1 _4936_ (.A(_3130_),
    .B(_3134_),
    .C(_0966_),
    .D(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__buf_6 _4937_ (.A(_0873_),
    .X(_0972_));
 sky130_fd_sc_hd__o221ai_4 _4938_ (.A1(_0964_),
    .A2(_0965_),
    .B1(_0971_),
    .B2(_3126_),
    .C1(net17),
    .Y(_0973_));
 sky130_fd_sc_hd__or3_2 _4939_ (.A(_0873_),
    .B(_0964_),
    .C(_0965_),
    .X(_0974_));
 sky130_fd_sc_hd__and2_0 _4940_ (.A(_0973_),
    .B(_0974_),
    .X(_2982_));
 sky130_fd_sc_hd__o21ai_0 _4941_ (.A1(_2811_),
    .A2(_0887_),
    .B1(_2808_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2b_2 _4942_ (.A_N(_2807_),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__xor2_4 _4943_ (.A(_2942_),
    .B(_0976_),
    .X(_3029_));
 sky130_fd_sc_hd__or2_1 _4944_ (.A(_0964_),
    .B(_0965_),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _4945_ (.A(_3134_),
    .B(_0970_),
    .Y(_0978_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_3025_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__nor3_1 _4947_ (.A(_3126_),
    .B(_3130_),
    .C(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _4948_ (.A(_3057_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__a21boi_0 _4949_ (.A1(_0977_),
    .A2(_0981_),
    .B1_N(_0974_),
    .Y(_3030_));
 sky130_fd_sc_hd__and2_0 _4950_ (.A(_0973_),
    .B(_0974_),
    .X(_3033_));
 sky130_fd_sc_hd__xor2_1 _4951_ (.A(_0977_),
    .B(_0981_),
    .X(_2985_));
 sky130_fd_sc_hd__buf_6 _4952_ (.A(_0972_),
    .X(_3038_));
 sky130_fd_sc_hd__nand2_1 _4953_ (.A(net24),
    .B(_0971_),
    .Y(_0982_));
 sky130_fd_sc_hd__xor2_1 _4954_ (.A(_3126_),
    .B(_0982_),
    .X(_2991_));
 sky130_fd_sc_hd__nand2_1 _4955_ (.A(net24),
    .B(_0979_),
    .Y(_0983_));
 sky130_fd_sc_hd__xor2_1 _4956_ (.A(_3130_),
    .B(_0983_),
    .X(_2995_));
 sky130_fd_sc_hd__o21ai_0 _4957_ (.A1(_0966_),
    .A2(_0970_),
    .B1(net17),
    .Y(_0984_));
 sky130_fd_sc_hd__xor2_1 _4958_ (.A(_3134_),
    .B(_0984_),
    .X(_2999_));
 sky130_fd_sc_hd__a21oi_1 _4959_ (.A1(_3025_),
    .A2(_0969_),
    .B1(_3057_),
    .Y(_0985_));
 sky130_fd_sc_hd__xnor2_1 _4960_ (.A(_3152_),
    .B(_0985_),
    .Y(_3003_));
 sky130_fd_sc_hd__o21ai_0 _4961_ (.A1(_0966_),
    .A2(_0968_),
    .B1(net17),
    .Y(_0986_));
 sky130_fd_sc_hd__xor2_1 _4962_ (.A(_3138_),
    .B(_0986_),
    .X(_3007_));
 sky130_fd_sc_hd__a21oi_1 _4963_ (.A1(_3025_),
    .A2(_0967_),
    .B1(_3057_),
    .Y(_0987_));
 sky130_fd_sc_hd__xnor2_1 _4964_ (.A(_3142_),
    .B(_0987_),
    .Y(_3011_));
 sky130_fd_sc_hd__o21ai_0 _4965_ (.A1(_0966_),
    .A2(_3082_),
    .B1(_0972_),
    .Y(_0988_));
 sky130_fd_sc_hd__xor2_1 _4966_ (.A(_3146_),
    .B(_0988_),
    .X(_3015_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_3025_),
    .B(_3057_),
    .Y(_0989_));
 sky130_fd_sc_hd__xnor2_1 _4968_ (.A(_3082_),
    .B(_0989_),
    .Y(_3019_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_3026_),
    .B(net26),
    .Y(_0990_));
 sky130_fd_sc_hd__o21ai_2 _4970_ (.A1(_0972_),
    .A2(_3023_),
    .B1(_0990_),
    .Y(_2151_));
 sky130_fd_sc_hd__inv_1 _4971_ (.A(_2151_),
    .Y(_2155_));
 sky130_fd_sc_hd__inv_1 _4972_ (.A(_3021_),
    .Y(_0991_));
 sky130_fd_sc_hd__nor2b_1 _4973_ (.A(_2150_),
    .B_N(_3028_),
    .Y(_0992_));
 sky130_fd_sc_hd__o21ai_0 _4974_ (.A1(_3027_),
    .A2(_0992_),
    .B1(_3022_),
    .Y(_0993_));
 sky130_fd_sc_hd__a21boi_0 _4975_ (.A1(_0991_),
    .A2(_0993_),
    .B1_N(_3018_),
    .Y(_0994_));
 sky130_fd_sc_hd__o21ai_0 _4976_ (.A1(_3017_),
    .A2(_0994_),
    .B1(_3014_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2b_1 _4977_ (.A_N(_3013_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__a21o_1 _4978_ (.A1(_3010_),
    .A2(_0996_),
    .B1(_3009_),
    .X(_0997_));
 sky130_fd_sc_hd__a21o_1 _4979_ (.A1(_3006_),
    .A2(_0997_),
    .B1(_3005_),
    .X(_0998_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_3002_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2b_1 _4981_ (.A_N(_3001_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a21o_1 _4982_ (.A1(_2998_),
    .A2(_1000_),
    .B1(_2997_),
    .X(_1001_));
 sky130_fd_sc_hd__nand3_1 _4983_ (.A(_2990_),
    .B(_2994_),
    .C(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__a21oi_1 _4984_ (.A1(_2988_),
    .A2(_2993_),
    .B1(_2987_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__a21o_1 _4986_ (.A1(_3036_),
    .A2(_1004_),
    .B1(_3035_),
    .X(_1005_));
 sky130_fd_sc_hd__a21oi_1 _4987_ (.A1(_3032_),
    .A2(_1005_),
    .B1(_3031_),
    .Y(_1006_));
 sky130_fd_sc_hd__xnor2_2 _4988_ (.A(_2984_),
    .B(_1006_),
    .Y(_3197_));
 sky130_fd_sc_hd__inv_1 _4989_ (.A(_2993_),
    .Y(_1007_));
 sky130_fd_sc_hd__nor2b_1 _4990_ (.A(_2152_),
    .B_N(_3022_),
    .Y(_1008_));
 sky130_fd_sc_hd__o21ai_0 _4991_ (.A1(_3021_),
    .A2(_1008_),
    .B1(_3018_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2b_1 _4992_ (.A_N(_3017_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__a21o_1 _4993_ (.A1(_3014_),
    .A2(_1010_),
    .B1(_3013_),
    .X(_1011_));
 sky130_fd_sc_hd__a21o_1 _4994_ (.A1(_3010_),
    .A2(_1011_),
    .B1(_3009_),
    .X(_1012_));
 sky130_fd_sc_hd__a21o_1 _4995_ (.A1(_3006_),
    .A2(_1012_),
    .B1(_3005_),
    .X(_1013_));
 sky130_fd_sc_hd__a21o_1 _4996_ (.A1(_3002_),
    .A2(_1013_),
    .B1(_3001_),
    .X(_1014_));
 sky130_fd_sc_hd__a21o_1 _4997_ (.A1(_2998_),
    .A2(_1014_),
    .B1(_2997_),
    .X(_1015_));
 sky130_fd_sc_hd__nand2_1 _4998_ (.A(_2994_),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a21boi_1 _4999_ (.A1(_1007_),
    .A2(_1016_),
    .B1_N(_2990_),
    .Y(_1017_));
 sky130_fd_sc_hd__o21a_1 _5000_ (.A1(_2987_),
    .A2(_1017_),
    .B1(_3036_),
    .X(_1018_));
 sky130_fd_sc_hd__nor2_1 _5001_ (.A(_3035_),
    .B(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__xnor2_2 _5002_ (.A(_3032_),
    .B(_1019_),
    .Y(_3201_));
 sky130_fd_sc_hd__nand3_1 _5003_ (.A(_2998_),
    .B(_2990_),
    .C(_2994_),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_2 _5004_ (.A(_2994_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21oi_1 _5005_ (.A1(_2998_),
    .A2(_3001_),
    .B1(_2997_),
    .Y(_1022_));
 sky130_fd_sc_hd__o21ai_0 _5006_ (.A1(_1021_),
    .A2(_1022_),
    .B1(_1007_),
    .Y(_1023_));
 sky130_fd_sc_hd__a21oi_1 _5007_ (.A1(_2988_),
    .A2(_1023_),
    .B1(_2987_),
    .Y(_1024_));
 sky130_fd_sc_hd__o21ai_2 _5008_ (.A1(_0999_),
    .A2(_1020_),
    .B1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__xor2_4 _5009_ (.A(_3036_),
    .B(_1025_),
    .X(_3205_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_1007_),
    .B(_1016_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(_2990_),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_2 _5012_ (.A(_1017_),
    .B(_1027_),
    .Y(_3159_));
 sky130_fd_sc_hd__xnor2_4 _5013_ (.A(_1021_),
    .B(_1001_),
    .Y(_3209_));
 sky130_fd_sc_hd__xor2_2 _5014_ (.A(_3002_),
    .B(_0998_),
    .X(_3167_));
 sky130_fd_sc_hd__inv_1 _5015_ (.A(_3167_),
    .Y(_3108_));
 sky130_fd_sc_hd__xor2_4 _5016_ (.A(_3006_),
    .B(_1012_),
    .X(_3172_));
 sky130_fd_sc_hd__inv_1 _5017_ (.A(_3172_),
    .Y(_3109_));
 sky130_fd_sc_hd__inv_1 _5018_ (.A(_3045_),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_1 _5019_ (.A(_3051_),
    .Y(_1029_));
 sky130_fd_sc_hd__inv_1 _5020_ (.A(_3058_),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_1 _5021_ (.A(_3064_),
    .Y(_1031_));
 sky130_fd_sc_hd__inv_1 _5022_ (.A(_3070_),
    .Y(_1032_));
 sky130_fd_sc_hd__inv_1 _5023_ (.A(_3076_),
    .Y(_1033_));
 sky130_fd_sc_hd__nor2b_1 _5024_ (.A(net62),
    .B_N(_3080_),
    .Y(_1034_));
 sky130_fd_sc_hd__o21ai_1 _5025_ (.A1(_1034_),
    .A2(_3079_),
    .B1(_3077_),
    .Y(_1035_));
 sky130_fd_sc_hd__a21boi_2 _5026_ (.A1(_1035_),
    .A2(_1033_),
    .B1_N(_3074_),
    .Y(_1036_));
 sky130_fd_sc_hd__o21ai_2 _5027_ (.A1(_1036_),
    .A2(_3073_),
    .B1(_3071_),
    .Y(_1037_));
 sky130_fd_sc_hd__a21boi_2 _5028_ (.A1(_1037_),
    .A2(_1032_),
    .B1_N(_3068_),
    .Y(_1038_));
 sky130_fd_sc_hd__o21ai_2 _5029_ (.A1(_1038_),
    .A2(_3067_),
    .B1(_3065_),
    .Y(_1039_));
 sky130_fd_sc_hd__a21boi_2 _5030_ (.A1(_1039_),
    .A2(_1031_),
    .B1_N(_3062_),
    .Y(_1040_));
 sky130_fd_sc_hd__o21ai_2 _5031_ (.A1(_1040_),
    .A2(_3061_),
    .B1(_3059_),
    .Y(_1041_));
 sky130_fd_sc_hd__a21boi_2 _5032_ (.A1(_1041_),
    .A2(_1030_),
    .B1_N(_3055_),
    .Y(_1042_));
 sky130_fd_sc_hd__o21ai_2 _5033_ (.A1(_1042_),
    .A2(_3054_),
    .B1(_3052_),
    .Y(_1043_));
 sky130_fd_sc_hd__a21boi_2 _5034_ (.A1(_1043_),
    .A2(_1029_),
    .B1_N(_3049_),
    .Y(_1044_));
 sky130_fd_sc_hd__o21ai_2 _5035_ (.A1(_1044_),
    .A2(_3048_),
    .B1(_3046_),
    .Y(_1045_));
 sky130_fd_sc_hd__a21boi_2 _5036_ (.A1(_1028_),
    .A2(_1045_),
    .B1_N(_3043_),
    .Y(_1046_));
 sky130_fd_sc_hd__o21a_1 _5037_ (.A1(_3042_),
    .A2(_1046_),
    .B1(_3040_),
    .X(_1047_));
 sky130_fd_sc_hd__or2_4 _5038_ (.A(_3039_),
    .B(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__buf_12 _5039_ (.A(_1048_),
    .X(_3213_));
 sky130_fd_sc_hd__clkinv_8 _5040_ (.A(_3213_),
    .Y(_1049_));
 sky130_fd_sc_hd__buf_12 _5041_ (.A(_1049_),
    .X(_3235_));
 sky130_fd_sc_hd__inv_1 _5042_ (.A(_2905_),
    .Y(_1050_));
 sky130_fd_sc_hd__a21o_1 _5043_ (.A1(_2146_),
    .A2(_2923_),
    .B1(_2922_),
    .X(_1051_));
 sky130_fd_sc_hd__a21oi_1 _5044_ (.A1(_2917_),
    .A2(_1051_),
    .B1(_2916_),
    .Y(_1052_));
 sky130_fd_sc_hd__o21bai_1 _5045_ (.A1(_0891_),
    .A2(_1052_),
    .B1_N(_2912_),
    .Y(_1053_));
 sky130_fd_sc_hd__a21oi_1 _5046_ (.A1(_2909_),
    .A2(_1053_),
    .B1(_2908_),
    .Y(_1054_));
 sky130_fd_sc_hd__o21bai_1 _5047_ (.A1(_1050_),
    .A2(_1054_),
    .B1_N(_2904_),
    .Y(_1055_));
 sky130_fd_sc_hd__a21oi_2 _5048_ (.A1(_2902_),
    .A2(_1055_),
    .B1(_2901_),
    .Y(_1056_));
 sky130_fd_sc_hd__xnor2_2 _5049_ (.A(_3084_),
    .B(_1056_),
    .Y(_3086_));
 sky130_fd_sc_hd__inv_1 _5050_ (.A(_3086_),
    .Y(_3191_));
 sky130_fd_sc_hd__xor2_4 _5051_ (.A(_2998_),
    .B(_1014_),
    .X(_3163_));
 sky130_fd_sc_hd__inv_1 _5052_ (.A(_3095_),
    .Y(_1057_));
 sky130_fd_sc_hd__inv_1 _5053_ (.A(_3103_),
    .Y(_1058_));
 sky130_fd_sc_hd__a21o_1 _5054_ (.A1(_2156_),
    .A2(_3113_),
    .B1(_3112_),
    .X(_1059_));
 sky130_fd_sc_hd__a21oi_1 _5055_ (.A1(_3107_),
    .A2(_1059_),
    .B1(_3106_),
    .Y(_1060_));
 sky130_fd_sc_hd__o21bai_1 _5056_ (.A1(_1058_),
    .A2(_1060_),
    .B1_N(_3102_),
    .Y(_1061_));
 sky130_fd_sc_hd__a21oi_1 _5057_ (.A1(_3099_),
    .A2(_1061_),
    .B1(_3098_),
    .Y(_1062_));
 sky130_fd_sc_hd__o21bai_1 _5058_ (.A1(_1057_),
    .A2(_1062_),
    .B1_N(_3094_),
    .Y(_1063_));
 sky130_fd_sc_hd__a21oi_2 _5059_ (.A1(_3091_),
    .A2(_1063_),
    .B1(_3090_),
    .Y(_1064_));
 sky130_fd_sc_hd__xnor2_2 _5060_ (.A(_3088_),
    .B(_1064_),
    .Y(_3115_));
 sky130_fd_sc_hd__and2_0 _5061_ (.A(_0910_),
    .B(_0915_),
    .X(_3118_));
 sky130_fd_sc_hd__a21o_1 _5062_ (.A1(_2942_),
    .A2(_0976_),
    .B1(_2941_),
    .X(_1065_));
 sky130_fd_sc_hd__a21o_1 _5063_ (.A1(_2938_),
    .A2(_1065_),
    .B1(_2937_),
    .X(_1066_));
 sky130_fd_sc_hd__xor2_4 _5064_ (.A(_3120_),
    .B(_1066_),
    .X(_3121_));
 sky130_fd_sc_hd__a21boi_0 _5065_ (.A1(_0977_),
    .A2(_0981_),
    .B1_N(_0974_),
    .Y(_3122_));
 sky130_fd_sc_hd__inv_1 _5066_ (.A(_3150_),
    .Y(_1067_));
 sky130_fd_sc_hd__inv_1 _5067_ (.A(_3140_),
    .Y(_1068_));
 sky130_fd_sc_hd__inv_1 _5068_ (.A(_3148_),
    .Y(_1069_));
 sky130_fd_sc_hd__inv_1 _5069_ (.A(_2902_),
    .Y(_1070_));
 sky130_fd_sc_hd__o21bai_1 _5070_ (.A1(_1070_),
    .A2(_0896_),
    .B1_N(_2901_),
    .Y(_1071_));
 sky130_fd_sc_hd__a21oi_1 _5071_ (.A1(_3084_),
    .A2(_1071_),
    .B1(_3083_),
    .Y(_1072_));
 sky130_fd_sc_hd__o21bai_1 _5072_ (.A1(_1069_),
    .A2(_1072_),
    .B1_N(_3147_),
    .Y(_1073_));
 sky130_fd_sc_hd__a21oi_1 _5073_ (.A1(_3144_),
    .A2(_1073_),
    .B1(_3143_),
    .Y(_1074_));
 sky130_fd_sc_hd__o21bai_1 _5074_ (.A1(_1068_),
    .A2(_1074_),
    .B1_N(_3139_),
    .Y(_1075_));
 sky130_fd_sc_hd__a21oi_2 _5075_ (.A1(_3154_),
    .A2(_1075_),
    .B1(_3153_),
    .Y(_1076_));
 sky130_fd_sc_hd__o21bai_1 _5076_ (.A1(_1067_),
    .A2(_1076_),
    .B1_N(_3135_),
    .Y(_1077_));
 sky130_fd_sc_hd__a21oi_2 _5077_ (.A1(_3132_),
    .A2(_1077_),
    .B1(_3131_),
    .Y(_1078_));
 sky130_fd_sc_hd__xnor2_4 _5078_ (.A(_3128_),
    .B(_1078_),
    .Y(_3294_));
 sky130_fd_sc_hd__inv_1 _5079_ (.A(_3132_),
    .Y(_1079_));
 sky130_fd_sc_hd__inv_1 _5080_ (.A(_3154_),
    .Y(_1080_));
 sky130_fd_sc_hd__inv_1 _5081_ (.A(_3144_),
    .Y(_1081_));
 sky130_fd_sc_hd__inv_1 _5082_ (.A(_3084_),
    .Y(_1082_));
 sky130_fd_sc_hd__o21bai_1 _5083_ (.A1(_1082_),
    .A2(_1056_),
    .B1_N(_3083_),
    .Y(_1083_));
 sky130_fd_sc_hd__a21oi_2 _5084_ (.A1(_3148_),
    .A2(_1083_),
    .B1(_3147_),
    .Y(_1084_));
 sky130_fd_sc_hd__o21bai_1 _5085_ (.A1(_1081_),
    .A2(_1084_),
    .B1_N(_3143_),
    .Y(_1085_));
 sky130_fd_sc_hd__a21oi_2 _5086_ (.A1(_3140_),
    .A2(_1085_),
    .B1(_3139_),
    .Y(_1086_));
 sky130_fd_sc_hd__o21bai_1 _5087_ (.A1(_1080_),
    .A2(_1086_),
    .B1_N(_3153_),
    .Y(_1087_));
 sky130_fd_sc_hd__a21oi_2 _5088_ (.A1(_3136_),
    .A2(_1087_),
    .B1(_3135_),
    .Y(_1088_));
 sky130_fd_sc_hd__xnor2_2 _5089_ (.A(_1079_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__inv_1 _5090_ (.A(_1089_),
    .Y(_3310_));
 sky130_fd_sc_hd__xnor2_4 _5091_ (.A(_3150_),
    .B(_1076_),
    .Y(_3298_));
 sky130_fd_sc_hd__xnor2_2 _5092_ (.A(_3154_),
    .B(_1086_),
    .Y(_3316_));
 sky130_fd_sc_hd__xnor2_2 _5093_ (.A(_3140_),
    .B(_1074_),
    .Y(_3302_));
 sky130_fd_sc_hd__xnor2_2 _5094_ (.A(_3144_),
    .B(_1084_),
    .Y(_3306_));
 sky130_fd_sc_hd__inv_1 _5095_ (.A(_3032_),
    .Y(_1090_));
 sky130_fd_sc_hd__o21bai_1 _5096_ (.A1(_1090_),
    .A2(_1019_),
    .B1_N(_3031_),
    .Y(_1091_));
 sky130_fd_sc_hd__a21o_1 _5097_ (.A1(_2984_),
    .A2(_1091_),
    .B1(_2983_),
    .X(_1092_));
 sky130_fd_sc_hd__xor2_1 _5098_ (.A(_3124_),
    .B(_1092_),
    .X(_3156_));
 sky130_fd_sc_hd__xnor2_2 _5099_ (.A(_3148_),
    .B(_1072_),
    .Y(_3257_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_2938_),
    .B(_3120_),
    .Y(_1093_));
 sky130_fd_sc_hd__a21oi_1 _5101_ (.A1(_3120_),
    .A2(_2937_),
    .B1(_3119_),
    .Y(_1094_));
 sky130_fd_sc_hd__o21ai_0 _5102_ (.A1(_0917_),
    .A2(_1093_),
    .B1(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__o21ba_1 _5103_ (.A1(_0950_),
    .A2(_0951_),
    .B1_N(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nor3b_2 _5104_ (.A(_0950_),
    .B(_0951_),
    .C_N(_1095_),
    .Y(_1097_));
 sky130_fd_sc_hd__a211oi_2 _5105_ (.A1(_0909_),
    .A2(_0910_),
    .B1(_1096_),
    .C1(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__o211a_1 _5106_ (.A1(_1096_),
    .A2(_1097_),
    .B1(_0909_),
    .C1(_0910_),
    .X(_1099_));
 sky130_fd_sc_hd__nor3_1 _5107_ (.A(_3000_),
    .B(_3004_),
    .C(_3008_),
    .Y(_1100_));
 sky130_fd_sc_hd__inv_1 _5108_ (.A(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__or2_0 _5109_ (.A(_2992_),
    .B(_2996_),
    .X(_1102_));
 sky130_fd_sc_hd__or4_1 _5110_ (.A(_3034_),
    .B(_2986_),
    .C(_1101_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__o41ai_1 _5111_ (.A1(_2981_),
    .A2(_3029_),
    .A3(_3121_),
    .A4(_1103_),
    .B1(net17),
    .Y(_1104_));
 sky130_fd_sc_hd__nor3_2 _5112_ (.A(_1098_),
    .B(_1099_),
    .C(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__o21a_2 _5113_ (.A1(_1098_),
    .A2(_1099_),
    .B1(_3057_),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_0952_),
    .B(_0958_),
    .Y(_2973_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_0962_),
    .B(_0963_),
    .Y(_1107_));
 sky130_fd_sc_hd__o21bai_1 _5116_ (.A1(_1079_),
    .A2(_1088_),
    .B1_N(_3131_),
    .Y(_1108_));
 sky130_fd_sc_hd__a21oi_2 _5117_ (.A1(_3128_),
    .A2(_1108_),
    .B1(_3127_),
    .Y(_1109_));
 sky130_fd_sc_hd__xnor3_4 _5118_ (.A(_2973_),
    .B(_1107_),
    .C(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__o21a_1 _5119_ (.A1(_1105_),
    .A2(_1106_),
    .B1(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__nor3_4 _5120_ (.A(_1105_),
    .B(_1106_),
    .C(_1110_),
    .Y(_1112_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(_1111_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__nor2_1 _5122_ (.A(_3306_),
    .B(_3257_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2_1 _5123_ (.A(_3193_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__nor3_1 _5124_ (.A(_3316_),
    .B(_3302_),
    .C(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__nor2b_1 _5125_ (.A(_3298_),
    .B_N(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a21oi_1 _5126_ (.A1(_1089_),
    .A2(_1117_),
    .B1(net25),
    .Y(_1118_));
 sky130_fd_sc_hd__nor2_1 _5127_ (.A(_3294_),
    .B(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_1 _5128_ (.A(net11),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor3_4 _5129_ (.A(_1111_),
    .B(net10),
    .C(_1112_),
    .Y(_1121_));
 sky130_fd_sc_hd__a21oi_1 _5130_ (.A1(_1113_),
    .A2(_1120_),
    .B1(_1121_),
    .Y(_3155_));
 sky130_fd_sc_hd__inv_1 _5131_ (.A(_3302_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand4_1 _5132_ (.A(_3192_),
    .B(_3191_),
    .C(_1122_),
    .D(_1114_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor3_1 _5133_ (.A(_3298_),
    .B(_3316_),
    .C(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_1089_),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__nor2_1 _5135_ (.A(_3294_),
    .B(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__nor2_1 _5136_ (.A(net25),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__o21a_2 _5137_ (.A1(_1111_),
    .A2(_1112_),
    .B1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__nor2_2 _5138_ (.A(_1121_),
    .B(_1128_),
    .Y(_3198_));
 sky130_fd_sc_hd__a21oi_1 _5139_ (.A1(_1113_),
    .A2(_1120_),
    .B1(_1121_),
    .Y(_3202_));
 sky130_fd_sc_hd__nor2_1 _5140_ (.A(_1121_),
    .B(_1128_),
    .Y(_3206_));
 sky130_fd_sc_hd__a21oi_1 _5141_ (.A1(_1113_),
    .A2(_1120_),
    .B1(_1121_),
    .Y(_3160_));
 sky130_fd_sc_hd__nor2_1 _5142_ (.A(_1113_),
    .B(_1127_),
    .Y(_1129_));
 sky130_fd_sc_hd__nor2_1 _5143_ (.A(_1128_),
    .B(_1129_),
    .Y(_3210_));
 sky130_fd_sc_hd__xnor2_1 _5144_ (.A(_3294_),
    .B(_1118_),
    .Y(_3164_));
 sky130_fd_sc_hd__nor2_1 _5145_ (.A(net11),
    .B(_1124_),
    .Y(_1130_));
 sky130_fd_sc_hd__xnor2_1 _5146_ (.A(_3310_),
    .B(_1130_),
    .Y(_3168_));
 sky130_fd_sc_hd__nor2_1 _5147_ (.A(net11),
    .B(_1116_),
    .Y(_1131_));
 sky130_fd_sc_hd__xnor2_1 _5148_ (.A(_3298_),
    .B(_1131_),
    .Y(_3171_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(net10),
    .B(_1123_),
    .Y(_1132_));
 sky130_fd_sc_hd__xor2_1 _5150_ (.A(_3316_),
    .B(_1132_),
    .X(_3175_));
 sky130_fd_sc_hd__nand2_1 _5151_ (.A(net19),
    .B(_1115_),
    .Y(_1133_));
 sky130_fd_sc_hd__xnor2_1 _5152_ (.A(_1122_),
    .B(_1133_),
    .Y(_3179_));
 sky130_fd_sc_hd__nor3_1 _5153_ (.A(_2925_),
    .B(_3086_),
    .C(_3257_),
    .Y(_1134_));
 sky130_fd_sc_hd__nor2_1 _5154_ (.A(net11),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__xnor2_1 _5155_ (.A(_3306_),
    .B(_1135_),
    .Y(_3184_));
 sky130_fd_sc_hd__nor2_1 _5156_ (.A(_3193_),
    .B(_3235_),
    .Y(_1136_));
 sky130_fd_sc_hd__xnor2_1 _5157_ (.A(_3257_),
    .B(_1136_),
    .Y(_3187_));
 sky130_fd_sc_hd__mux2i_4 _5158_ (.A0(_3194_),
    .A1(_3086_),
    .S(_3235_),
    .Y(_2161_));
 sky130_fd_sc_hd__inv_1 _5159_ (.A(_3204_),
    .Y(_1137_));
 sky130_fd_sc_hd__inv_1 _5160_ (.A(_3162_),
    .Y(_1138_));
 sky130_fd_sc_hd__inv_1 _5161_ (.A(_3166_),
    .Y(_1139_));
 sky130_fd_sc_hd__inv_1 _5162_ (.A(_3174_),
    .Y(_1140_));
 sky130_fd_sc_hd__inv_1 _5163_ (.A(_3182_),
    .Y(_1141_));
 sky130_fd_sc_hd__a21o_1 _5164_ (.A1(_2163_),
    .A2(_3190_),
    .B1(_3189_),
    .X(_1142_));
 sky130_fd_sc_hd__a21oi_1 _5165_ (.A1(_3186_),
    .A2(_1142_),
    .B1(_3185_),
    .Y(_1143_));
 sky130_fd_sc_hd__o21bai_1 _5166_ (.A1(_1141_),
    .A2(_1143_),
    .B1_N(_3181_),
    .Y(_1144_));
 sky130_fd_sc_hd__a21oi_1 _5167_ (.A1(_3178_),
    .A2(_1144_),
    .B1(_3177_),
    .Y(_1145_));
 sky130_fd_sc_hd__o21bai_1 _5168_ (.A1(_1140_),
    .A2(_1145_),
    .B1_N(_3173_),
    .Y(_1146_));
 sky130_fd_sc_hd__a21oi_2 _5169_ (.A1(_3170_),
    .A2(_1146_),
    .B1(_3169_),
    .Y(_1147_));
 sky130_fd_sc_hd__o21bai_1 _5170_ (.A1(_1139_),
    .A2(_1147_),
    .B1_N(_3165_),
    .Y(_1148_));
 sky130_fd_sc_hd__a21oi_2 _5171_ (.A1(_3212_),
    .A2(_1148_),
    .B1(_3211_),
    .Y(_1149_));
 sky130_fd_sc_hd__o21bai_1 _5172_ (.A1(_1138_),
    .A2(_1149_),
    .B1_N(_3161_),
    .Y(_1150_));
 sky130_fd_sc_hd__a21oi_2 _5173_ (.A1(_3208_),
    .A2(_1150_),
    .B1(_3207_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21bai_1 _5174_ (.A1(_1137_),
    .A2(_1151_),
    .B1_N(_3203_),
    .Y(_1152_));
 sky130_fd_sc_hd__a21oi_2 _5175_ (.A1(_3200_),
    .A2(_1152_),
    .B1(_3199_),
    .Y(_1153_));
 sky130_fd_sc_hd__xnor2_4 _5176_ (.A(_3158_),
    .B(_1153_),
    .Y(_3321_));
 sky130_fd_sc_hd__inv_1 _5177_ (.A(_2165_),
    .Y(_2162_));
 sky130_fd_sc_hd__a21o_1 _5178_ (.A1(_2162_),
    .A2(_3196_),
    .B1(_3195_),
    .X(_1154_));
 sky130_fd_sc_hd__a21o_1 _5179_ (.A1(_3190_),
    .A2(_1154_),
    .B1(_3189_),
    .X(_1155_));
 sky130_fd_sc_hd__a21oi_2 _5180_ (.A1(_1155_),
    .A2(_3186_),
    .B1(_3185_),
    .Y(_1156_));
 sky130_fd_sc_hd__o21bai_2 _5181_ (.A1(_1141_),
    .A2(_1156_),
    .B1_N(_3181_),
    .Y(_1157_));
 sky130_fd_sc_hd__a21oi_2 _5182_ (.A1(_3178_),
    .A2(_1157_),
    .B1(_3177_),
    .Y(_1158_));
 sky130_fd_sc_hd__o21bai_2 _5183_ (.A1(_1140_),
    .A2(_1158_),
    .B1_N(_3173_),
    .Y(_1159_));
 sky130_fd_sc_hd__a21oi_2 _5184_ (.A1(_1159_),
    .A2(_3170_),
    .B1(_3169_),
    .Y(_1160_));
 sky130_fd_sc_hd__o21bai_4 _5185_ (.A1(_1139_),
    .A2(_1160_),
    .B1_N(_3165_),
    .Y(_1161_));
 sky130_fd_sc_hd__a21oi_2 _5186_ (.A1(_1161_),
    .A2(_3212_),
    .B1(_3211_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21bai_4 _5187_ (.A1(_1138_),
    .A2(_1162_),
    .B1_N(_3161_),
    .Y(_1163_));
 sky130_fd_sc_hd__a21oi_2 _5188_ (.A1(_3208_),
    .A2(_1163_),
    .B1(_3207_),
    .Y(_1164_));
 sky130_fd_sc_hd__o21bai_4 _5189_ (.A1(_1164_),
    .A2(_1137_),
    .B1_N(_3203_),
    .Y(_1165_));
 sky130_fd_sc_hd__xor2_4 _5190_ (.A(_3200_),
    .B(_1165_),
    .X(_3361_));
 sky130_fd_sc_hd__xnor2_4 _5191_ (.A(_3204_),
    .B(_1151_),
    .Y(_3365_));
 sky130_fd_sc_hd__xor2_4 _5192_ (.A(_3208_),
    .B(_1163_),
    .X(_3368_));
 sky130_fd_sc_hd__xnor2_4 _5193_ (.A(_3162_),
    .B(_1149_),
    .Y(_3324_));
 sky130_fd_sc_hd__xor2_4 _5194_ (.A(_3212_),
    .B(_1161_),
    .X(_3372_));
 sky130_fd_sc_hd__xnor2_2 _5195_ (.A(_3166_),
    .B(_1147_),
    .Y(_3328_));
 sky130_fd_sc_hd__xor2_2 _5196_ (.A(_3170_),
    .B(_1159_),
    .X(_3376_));
 sky130_fd_sc_hd__inv_1 _5197_ (.A(_3219_),
    .Y(_1166_));
 sky130_fd_sc_hd__inv_1 _5198_ (.A(_3225_),
    .Y(_1167_));
 sky130_fd_sc_hd__inv_1 _5199_ (.A(_3231_),
    .Y(_1168_));
 sky130_fd_sc_hd__inv_1 _5200_ (.A(_3238_),
    .Y(_1169_));
 sky130_fd_sc_hd__inv_1 _5201_ (.A(_3244_),
    .Y(_1170_));
 sky130_fd_sc_hd__inv_1 _5202_ (.A(_3250_),
    .Y(_1171_));
 sky130_fd_sc_hd__a21o_1 _5203_ (.A1(_3256_),
    .A2(net62),
    .B1(_3255_),
    .X(_1172_));
 sky130_fd_sc_hd__a21oi_2 _5204_ (.A1(_1172_),
    .A2(_3253_),
    .B1(_3252_),
    .Y(_1173_));
 sky130_fd_sc_hd__o21bai_1 _5205_ (.A1(_1173_),
    .A2(_1171_),
    .B1_N(_3249_),
    .Y(_1174_));
 sky130_fd_sc_hd__a21oi_2 _5206_ (.A1(_1174_),
    .A2(_3247_),
    .B1(_3246_),
    .Y(_1175_));
 sky130_fd_sc_hd__o21bai_1 _5207_ (.A1(_1175_),
    .A2(_1170_),
    .B1_N(_3243_),
    .Y(_1176_));
 sky130_fd_sc_hd__a21oi_2 _5208_ (.A1(_1176_),
    .A2(_3241_),
    .B1(_3240_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21bai_1 _5209_ (.A1(_1177_),
    .A2(_1169_),
    .B1_N(_3237_),
    .Y(_1178_));
 sky130_fd_sc_hd__a21oi_2 _5210_ (.A1(_1178_),
    .A2(_3234_),
    .B1(_3233_),
    .Y(_1179_));
 sky130_fd_sc_hd__o21bai_1 _5211_ (.A1(_1179_),
    .A2(_1168_),
    .B1_N(_3230_),
    .Y(_1180_));
 sky130_fd_sc_hd__a21oi_2 _5212_ (.A1(_1180_),
    .A2(_3228_),
    .B1(_3227_),
    .Y(_1181_));
 sky130_fd_sc_hd__o21bai_1 _5213_ (.A1(_1167_),
    .A2(_1181_),
    .B1_N(_3224_),
    .Y(_1182_));
 sky130_fd_sc_hd__a21oi_2 _5214_ (.A1(_1182_),
    .A2(_3222_),
    .B1(_3221_),
    .Y(_1183_));
 sky130_fd_sc_hd__o21bai_1 _5215_ (.A1(_1183_),
    .A2(_1166_),
    .B1_N(_3218_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21o_2 _5216_ (.A1(_1184_),
    .A2(_3216_),
    .B1(_3215_),
    .X(_1185_));
 sky130_fd_sc_hd__inv_4 _5217_ (.A(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__buf_8 _5218_ (.A(_1186_),
    .X(_3405_));
 sky130_fd_sc_hd__inv_1 _5219_ (.A(_3091_),
    .Y(_1187_));
 sky130_fd_sc_hd__inv_1 _5220_ (.A(_3099_),
    .Y(_1188_));
 sky130_fd_sc_hd__a21oi_1 _5221_ (.A1(_3107_),
    .A2(_2158_),
    .B1(_3106_),
    .Y(_1189_));
 sky130_fd_sc_hd__nor2_1 _5222_ (.A(_1058_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _5223_ (.A(_3102_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o21bai_1 _5224_ (.A1(_1188_),
    .A2(_1191_),
    .B1_N(_3098_),
    .Y(_1192_));
 sky130_fd_sc_hd__a21oi_1 _5225_ (.A1(_3095_),
    .A2(_1192_),
    .B1(_3094_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21bai_1 _5226_ (.A1(_1187_),
    .A2(_1193_),
    .B1_N(_3090_),
    .Y(_1194_));
 sky130_fd_sc_hd__a21oi_2 _5227_ (.A1(_3088_),
    .A2(_1194_),
    .B1(_3087_),
    .Y(_1195_));
 sky130_fd_sc_hd__xnor2_2 _5228_ (.A(_3260_),
    .B(_1195_),
    .Y(_3262_));
 sky130_fd_sc_hd__inv_1 _5229_ (.A(_3376_),
    .Y(_3286_));
 sky130_fd_sc_hd__inv_1 _5230_ (.A(_3328_),
    .Y(_3285_));
 sky130_fd_sc_hd__inv_1 _5231_ (.A(_3268_),
    .Y(_1196_));
 sky130_fd_sc_hd__inv_1 _5232_ (.A(_3276_),
    .Y(_1197_));
 sky130_fd_sc_hd__inv_1 _5233_ (.A(_3280_),
    .Y(_1198_));
 sky130_fd_sc_hd__a21oi_1 _5234_ (.A1(_2168_),
    .A2(_3284_),
    .B1(_3283_),
    .Y(_1199_));
 sky130_fd_sc_hd__nor2_1 _5235_ (.A(_1198_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nor2_1 _5236_ (.A(_3279_),
    .B(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__o21bai_1 _5237_ (.A1(_1197_),
    .A2(_1201_),
    .B1_N(_3275_),
    .Y(_1202_));
 sky130_fd_sc_hd__a21oi_2 _5238_ (.A1(_3272_),
    .A2(_1202_),
    .B1(_3271_),
    .Y(_1203_));
 sky130_fd_sc_hd__o21bai_1 _5239_ (.A1(_1196_),
    .A2(_1203_),
    .B1_N(_3267_),
    .Y(_1204_));
 sky130_fd_sc_hd__a21oi_2 _5240_ (.A1(_1204_),
    .A2(_3432_),
    .B1(_3431_),
    .Y(_1205_));
 sky130_fd_sc_hd__xnor2_4 _5241_ (.A(net113),
    .B(net194),
    .Y(_3292_));
 sky130_fd_sc_hd__inv_1 _5242_ (.A(_3292_),
    .Y(_3460_));
 sky130_fd_sc_hd__inv_1 _5243_ (.A(_3315_),
    .Y(_1206_));
 sky130_fd_sc_hd__inv_1 _5244_ (.A(_3305_),
    .Y(_1207_));
 sky130_fd_sc_hd__inv_1 _5245_ (.A(_3260_),
    .Y(_1208_));
 sky130_fd_sc_hd__o21bai_1 _5246_ (.A1(_1208_),
    .A2(_1195_),
    .B1_N(_3259_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21oi_2 _5247_ (.A1(_3309_),
    .A2(_1209_),
    .B1(_3308_),
    .Y(_1210_));
 sky130_fd_sc_hd__o21bai_1 _5248_ (.A1(_1207_),
    .A2(_1210_),
    .B1_N(_3304_),
    .Y(_1211_));
 sky130_fd_sc_hd__a21oi_2 _5249_ (.A1(_3319_),
    .A2(_1211_),
    .B1(_3318_),
    .Y(_1212_));
 sky130_fd_sc_hd__o21bai_1 _5250_ (.A1(_1206_),
    .A2(_1212_),
    .B1_N(_3300_),
    .Y(_1213_));
 sky130_fd_sc_hd__a21oi_2 _5251_ (.A1(_3313_),
    .A2(_1213_),
    .B1(_3312_),
    .Y(_1214_));
 sky130_fd_sc_hd__xnor2_4 _5252_ (.A(_3297_),
    .B(_1214_),
    .Y(_3581_));
 sky130_fd_sc_hd__inv_1 _5253_ (.A(_3319_),
    .Y(_1215_));
 sky130_fd_sc_hd__inv_1 _5254_ (.A(_3309_),
    .Y(_1216_));
 sky130_fd_sc_hd__inv_1 _5255_ (.A(_3088_),
    .Y(_1217_));
 sky130_fd_sc_hd__o21bai_1 _5256_ (.A1(_1217_),
    .A2(_1064_),
    .B1_N(_3087_),
    .Y(_1218_));
 sky130_fd_sc_hd__a21oi_2 _5257_ (.A1(_3260_),
    .A2(_1218_),
    .B1(_3259_),
    .Y(_1219_));
 sky130_fd_sc_hd__o21bai_1 _5258_ (.A1(_1216_),
    .A2(_1219_),
    .B1_N(_3308_),
    .Y(_1220_));
 sky130_fd_sc_hd__a21oi_2 _5259_ (.A1(_1220_),
    .A2(_3305_),
    .B1(_3304_),
    .Y(_1221_));
 sky130_fd_sc_hd__o21bai_1 _5260_ (.A1(_1215_),
    .A2(_1221_),
    .B1_N(_3318_),
    .Y(_1222_));
 sky130_fd_sc_hd__a21oi_2 _5261_ (.A1(_1222_),
    .A2(_3301_),
    .B1(_3300_),
    .Y(_1223_));
 sky130_fd_sc_hd__xnor2_4 _5262_ (.A(_3313_),
    .B(net114),
    .Y(_3565_));
 sky130_fd_sc_hd__xnor2_4 _5263_ (.A(_3315_),
    .B(_1212_),
    .Y(_3549_));
 sky130_fd_sc_hd__xnor2_4 _5264_ (.A(_3319_),
    .B(net128),
    .Y(_3533_));
 sky130_fd_sc_hd__xnor2_2 _5265_ (.A(_3305_),
    .B(_1210_),
    .Y(_3465_));
 sky130_fd_sc_hd__xnor2_2 _5266_ (.A(_3309_),
    .B(_1219_),
    .Y(_3424_));
 sky130_fd_sc_hd__inv_1 _5267_ (.A(_3115_),
    .Y(_3354_));
 sky130_fd_sc_hd__nor2_1 _5268_ (.A(_1096_),
    .B(_1097_),
    .Y(_1224_));
 sky130_fd_sc_hd__a21oi_1 _5269_ (.A1(_3036_),
    .A2(_1025_),
    .B1(_3035_),
    .Y(_1225_));
 sky130_fd_sc_hd__nor2_1 _5270_ (.A(_1090_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__o21ai_0 _5271_ (.A1(_3031_),
    .A2(_1226_),
    .B1(_2984_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand2b_1 _5272_ (.A_N(_2983_),
    .B(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__a21oi_1 _5273_ (.A1(_3124_),
    .A2(_1228_),
    .B1(_3123_),
    .Y(_1229_));
 sky130_fd_sc_hd__xnor3_4 _5274_ (.A(_2935_),
    .B(_1224_),
    .C(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__a21oi_2 _5275_ (.A1(_0973_),
    .A2(_0974_),
    .B1(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__and3_1 _5276_ (.A(_0973_),
    .B(_0974_),
    .C(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__nor3_4 _5277_ (.A(net10),
    .B(_1231_),
    .C(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__inv_1 _5278_ (.A(_3156_),
    .Y(_1234_));
 sky130_fd_sc_hd__nor3_2 _5279_ (.A(_3167_),
    .B(_3172_),
    .C(_3163_),
    .Y(_1235_));
 sky130_fd_sc_hd__nor3_1 _5280_ (.A(_3205_),
    .B(_3159_),
    .C(_3209_),
    .Y(_1236_));
 sky130_fd_sc_hd__nor2b_1 _5281_ (.A(_3201_),
    .B_N(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__nor2b_1 _5282_ (.A(_3197_),
    .B_N(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__a31oi_2 _5283_ (.A1(_1234_),
    .A2(_1235_),
    .A3(_1238_),
    .B1(net25),
    .Y(_1239_));
 sky130_fd_sc_hd__o21a_1 _5284_ (.A1(_1231_),
    .A2(_1232_),
    .B1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__or2_1 _5285_ (.A(_1105_),
    .B(_1106_),
    .X(_3129_));
 sky130_fd_sc_hd__inv_1 _5286_ (.A(_3313_),
    .Y(_1241_));
 sky130_fd_sc_hd__o21bai_1 _5287_ (.A1(_1241_),
    .A2(_1223_),
    .B1_N(_3312_),
    .Y(_1242_));
 sky130_fd_sc_hd__a21oi_1 _5288_ (.A1(_3297_),
    .A2(_1242_),
    .B1(_3296_),
    .Y(_1243_));
 sky130_fd_sc_hd__xnor3_4 _5289_ (.A(_3129_),
    .B(_1110_),
    .C(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__o21a_1 _5290_ (.A1(_1233_),
    .A2(_1240_),
    .B1(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__nor3_2 _5291_ (.A(_1233_),
    .B(_1240_),
    .C(_1244_),
    .Y(_1246_));
 sky130_fd_sc_hd__or2_0 _5292_ (.A(_1245_),
    .B(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_2 _5293_ (.A(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__nor2_1 _5294_ (.A(_3465_),
    .B(_3424_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _5295_ (.A(_3356_),
    .B(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__nor3_1 _5296_ (.A(_3549_),
    .B(_3533_),
    .C(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__nor2_1 _5297_ (.A(_3581_),
    .B(_3565_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21oi_2 _5298_ (.A1(_1251_),
    .A2(_1252_),
    .B1(_1186_),
    .Y(_1253_));
 sky130_fd_sc_hd__buf_6 _5299_ (.A(_1185_),
    .X(_3380_));
 sky130_fd_sc_hd__nor2_2 _5300_ (.A(net7),
    .B(_1248_),
    .Y(_1254_));
 sky130_fd_sc_hd__a21oi_1 _5301_ (.A1(_1248_),
    .A2(_1253_),
    .B1(_1254_),
    .Y(_3320_));
 sky130_fd_sc_hd__or3_1 _5302_ (.A(_3115_),
    .B(_3262_),
    .C(_3424_),
    .X(_1255_));
 sky130_fd_sc_hd__nor3_1 _5303_ (.A(_3533_),
    .B(_3465_),
    .C(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__or3b_1 _5304_ (.A(_3565_),
    .B(_3549_),
    .C_N(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__nor2_1 _5305_ (.A(_3581_),
    .B(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__nor2_2 _5306_ (.A(_1186_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__a21oi_1 _5307_ (.A1(_1248_),
    .A2(_1259_),
    .B1(_1254_),
    .Y(_3360_));
 sky130_fd_sc_hd__a21oi_1 _5308_ (.A1(_1248_),
    .A2(_1253_),
    .B1(_1254_),
    .Y(_3364_));
 sky130_fd_sc_hd__a21oi_1 _5309_ (.A1(_1248_),
    .A2(_1259_),
    .B1(_1254_),
    .Y(_3369_));
 sky130_fd_sc_hd__a21oi_1 _5310_ (.A1(_1248_),
    .A2(_1253_),
    .B1(_1254_),
    .Y(_3325_));
 sky130_fd_sc_hd__a21oi_1 _5311_ (.A1(_1248_),
    .A2(_1259_),
    .B1(_1254_),
    .Y(_3373_));
 sky130_fd_sc_hd__xor2_1 _5312_ (.A(_1248_),
    .B(_1253_),
    .X(_3329_));
 sky130_fd_sc_hd__nand2_1 _5313_ (.A(net20),
    .B(_1257_),
    .Y(_1260_));
 sky130_fd_sc_hd__xor2_1 _5314_ (.A(_3581_),
    .B(_1260_),
    .X(_3377_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_3405_),
    .B(_1251_),
    .Y(_1261_));
 sky130_fd_sc_hd__xnor2_1 _5316_ (.A(_3565_),
    .B(_1261_),
    .Y(_3333_));
 sky130_fd_sc_hd__nor2_1 _5317_ (.A(net8),
    .B(_1256_),
    .Y(_1262_));
 sky130_fd_sc_hd__xnor2_1 _5318_ (.A(_3549_),
    .B(_1262_),
    .Y(_3339_));
 sky130_fd_sc_hd__nand2_1 _5319_ (.A(net20),
    .B(_1250_),
    .Y(_1263_));
 sky130_fd_sc_hd__xor2_1 _5320_ (.A(_3533_),
    .B(_1263_),
    .X(_3342_));
 sky130_fd_sc_hd__nand2_1 _5321_ (.A(_3380_),
    .B(_1255_),
    .Y(_1264_));
 sky130_fd_sc_hd__xor2_1 _5322_ (.A(_3465_),
    .B(_1264_),
    .X(_3347_));
 sky130_fd_sc_hd__nor2_1 _5323_ (.A(_3356_),
    .B(_3405_),
    .Y(_1265_));
 sky130_fd_sc_hd__xnor2_1 _5324_ (.A(_3424_),
    .B(_1265_),
    .Y(_3351_));
 sky130_fd_sc_hd__inv_1 _5325_ (.A(_3262_),
    .Y(_3355_));
 sky130_fd_sc_hd__mux2i_4 _5326_ (.A0(_3357_),
    .A1(_3262_),
    .S(_3405_),
    .Y(_2171_));
 sky130_fd_sc_hd__inv_1 _5327_ (.A(_3367_),
    .Y(_1266_));
 sky130_fd_sc_hd__a21o_1 _5328_ (.A1(_2172_),
    .A2(_3353_),
    .B1(_3352_),
    .X(_1267_));
 sky130_fd_sc_hd__a21oi_2 _5329_ (.A1(_3349_),
    .A2(_1267_),
    .B1(_3348_),
    .Y(_1268_));
 sky130_fd_sc_hd__nor2b_1 _5330_ (.A(_1268_),
    .B_N(_3345_),
    .Y(_1269_));
 sky130_fd_sc_hd__o21ai_0 _5331_ (.A1(_3344_),
    .A2(_1269_),
    .B1(_3341_),
    .Y(_1270_));
 sky130_fd_sc_hd__nand2b_1 _5332_ (.A_N(_3340_),
    .B(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__a21o_1 _5333_ (.A1(_3337_),
    .A2(_1271_),
    .B1(_3334_),
    .X(_1272_));
 sky130_fd_sc_hd__a21oi_4 _5334_ (.A1(_3379_),
    .A2(_1272_),
    .B1(_3378_),
    .Y(_1273_));
 sky130_fd_sc_hd__nor2b_1 _5335_ (.A(_1273_),
    .B_N(_3331_),
    .Y(_1274_));
 sky130_fd_sc_hd__o21a_1 _5336_ (.A1(_3330_),
    .A2(_1274_),
    .B1(_3375_),
    .X(_1275_));
 sky130_fd_sc_hd__o21ai_0 _5337_ (.A1(_3374_),
    .A2(_1275_),
    .B1(_3327_),
    .Y(_1276_));
 sky130_fd_sc_hd__nand2b_1 _5338_ (.A_N(_3326_),
    .B(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__a21oi_2 _5339_ (.A1(_3371_),
    .A2(_1277_),
    .B1(_3370_),
    .Y(_1278_));
 sky130_fd_sc_hd__o21bai_1 _5340_ (.A1(_1266_),
    .A2(_1278_),
    .B1_N(_3366_),
    .Y(_1279_));
 sky130_fd_sc_hd__a21oi_2 _5341_ (.A1(_3363_),
    .A2(_1279_),
    .B1(_3362_),
    .Y(_1280_));
 sky130_fd_sc_hd__xnor2_2 _5342_ (.A(_3323_),
    .B(_1280_),
    .Y(_3665_));
 sky130_fd_sc_hd__inv_1 _5343_ (.A(_2174_),
    .Y(_2170_));
 sky130_fd_sc_hd__a21o_1 _5344_ (.A1(_3359_),
    .A2(_2170_),
    .B1(_3358_),
    .X(_1281_));
 sky130_fd_sc_hd__a21o_1 _5345_ (.A1(_1281_),
    .A2(_3353_),
    .B1(_3352_),
    .X(_1282_));
 sky130_fd_sc_hd__a21o_1 _5346_ (.A1(_3349_),
    .A2(_1282_),
    .B1(_3348_),
    .X(_1283_));
 sky130_fd_sc_hd__a21o_1 _5347_ (.A1(_1283_),
    .A2(_3345_),
    .B1(_3344_),
    .X(_1284_));
 sky130_fd_sc_hd__a21o_1 _5348_ (.A1(_3335_),
    .A2(_3340_),
    .B1(_3334_),
    .X(_1285_));
 sky130_fd_sc_hd__a31oi_4 _5349_ (.A1(_3341_),
    .A2(_1284_),
    .A3(_3337_),
    .B1(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__nor2b_1 _5350_ (.A(_1286_),
    .B_N(_3379_),
    .Y(_1287_));
 sky130_fd_sc_hd__o21ai_1 _5351_ (.A1(_1287_),
    .A2(_3378_),
    .B1(_3331_),
    .Y(_1288_));
 sky130_fd_sc_hd__nand2b_2 _5352_ (.A_N(_3330_),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__a21o_1 _5353_ (.A1(_1289_),
    .A2(_3375_),
    .B1(_3374_),
    .X(_1290_));
 sky130_fd_sc_hd__a21o_1 _5354_ (.A1(_1290_),
    .A2(_3327_),
    .B1(_3326_),
    .X(_1291_));
 sky130_fd_sc_hd__a21oi_2 _5355_ (.A1(_1291_),
    .A2(_3371_),
    .B1(_3370_),
    .Y(_1292_));
 sky130_fd_sc_hd__o21bai_2 _5356_ (.A1(_1266_),
    .A2(_1292_),
    .B1_N(_3366_),
    .Y(_1293_));
 sky130_fd_sc_hd__xor2_2 _5357_ (.A(_3363_),
    .B(net160),
    .X(_3657_));
 sky130_fd_sc_hd__xnor2_2 _5358_ (.A(_3367_),
    .B(_1278_),
    .Y(_3649_));
 sky130_fd_sc_hd__xor2_2 _5359_ (.A(_3371_),
    .B(net140),
    .X(_3641_));
 sky130_fd_sc_hd__nor2_1 _5360_ (.A(_3374_),
    .B(_1275_),
    .Y(_1294_));
 sky130_fd_sc_hd__xnor2_2 _5361_ (.A(_3327_),
    .B(_1294_),
    .Y(_3633_));
 sky130_fd_sc_hd__xnor2_4 _5362_ (.A(_3331_),
    .B(net264),
    .Y(_3620_));
 sky130_fd_sc_hd__inv_1 _5363_ (.A(_3389_),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_1 _5364_ (.A(_3400_),
    .Y(_1296_));
 sky130_fd_sc_hd__inv_1 _5365_ (.A(_3407_),
    .Y(_1297_));
 sky130_fd_sc_hd__inv_1 _5366_ (.A(_3413_),
    .Y(_1298_));
 sky130_fd_sc_hd__a21o_1 _5367_ (.A1(_3423_),
    .A2(_2122_),
    .B1(_3422_),
    .X(_1299_));
 sky130_fd_sc_hd__a21o_1 _5368_ (.A1(_1299_),
    .A2(_3420_),
    .B1(_3419_),
    .X(_1300_));
 sky130_fd_sc_hd__a21o_1 _5369_ (.A1(_1300_),
    .A2(_3417_),
    .B1(_3416_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_3414_),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__a21boi_2 _5371_ (.A1(_1302_),
    .A2(_1298_),
    .B1_N(_3411_),
    .Y(_1303_));
 sky130_fd_sc_hd__o21ai_1 _5372_ (.A1(_3410_),
    .A2(_1303_),
    .B1(_3408_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _5373_ (.A(_1304_),
    .B(_1297_),
    .Y(_1305_));
 sky130_fd_sc_hd__and2_4 _5374_ (.A(_1305_),
    .B(_3404_),
    .X(_1306_));
 sky130_fd_sc_hd__o21ai_2 _5375_ (.A1(_3403_),
    .A2(_1306_),
    .B1(_3401_),
    .Y(_1307_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(_1296_),
    .B(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__a21o_1 _5377_ (.A1(_1308_),
    .A2(_3398_),
    .B1(_3397_),
    .X(_1309_));
 sky130_fd_sc_hd__a21o_1 _5378_ (.A1(_1309_),
    .A2(_3395_),
    .B1(_3394_),
    .X(_1310_));
 sky130_fd_sc_hd__a21oi_2 _5379_ (.A1(_1310_),
    .A2(_3392_),
    .B1(_3391_),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_1 _5380_ (.A(_3388_),
    .Y(_1312_));
 sky130_fd_sc_hd__o21ai_2 _5381_ (.A1(_1295_),
    .A2(_1311_),
    .B1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a21o_1 _5382_ (.A1(_1313_),
    .A2(_3386_),
    .B1(_3385_),
    .X(_1314_));
 sky130_fd_sc_hd__nand2_2 _5383_ (.A(_1314_),
    .B(_3383_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2b_4 _5384_ (.A_N(_3382_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__buf_2 clone2 (.A(_0159_),
    .X(net2));
 sky130_fd_sc_hd__inv_8 _5386_ (.A(_1316_),
    .Y(_1318_));
 sky130_fd_sc_hd__buf_6 _5387_ (.A(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__buf_6 _5388_ (.A(_1319_),
    .X(_3517_));
 sky130_fd_sc_hd__or3_2 _5389_ (.A(net7),
    .B(_1245_),
    .C(_1246_),
    .X(_1320_));
 sky130_fd_sc_hd__o21ai_2 _5390_ (.A1(_1245_),
    .A2(_1246_),
    .B1(_1259_),
    .Y(_1321_));
 sky130_fd_sc_hd__a21o_1 _5391_ (.A1(_1165_),
    .A2(_3200_),
    .B1(_3199_),
    .X(_1322_));
 sky130_fd_sc_hd__a21oi_2 _5392_ (.A1(_1322_),
    .A2(_3158_),
    .B1(_3157_),
    .Y(_1323_));
 sky130_fd_sc_hd__xnor3_4 _5393_ (.A(_2982_),
    .B(_1230_),
    .C(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__a21o_1 _5394_ (.A1(_1293_),
    .A2(_3363_),
    .B1(_3362_),
    .X(_1325_));
 sky130_fd_sc_hd__a21oi_2 _5395_ (.A1(_1325_),
    .A2(_3323_),
    .B1(_3322_),
    .Y(_1326_));
 sky130_fd_sc_hd__xor3_2 _5396_ (.A(_3198_),
    .B(_1326_),
    .C(_1324_),
    .X(_1327_));
 sky130_fd_sc_hd__a21oi_4 _5397_ (.A1(_1320_),
    .A2(_1321_),
    .B1(net177),
    .Y(_1328_));
 sky130_fd_sc_hd__and3_4 _5398_ (.A(_1327_),
    .B(_1321_),
    .C(_1320_),
    .X(_1329_));
 sky130_fd_sc_hd__or2_4 _5399_ (.A(_1328_),
    .B(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__inv_4 _5400_ (.A(_1330_),
    .Y(_3441_));
 sky130_fd_sc_hd__inv_1 _5401_ (.A(_3272_),
    .Y(_1331_));
 sky130_fd_sc_hd__a21o_1 _5402_ (.A1(_2166_),
    .A2(_3290_),
    .B1(_3289_),
    .X(_1332_));
 sky130_fd_sc_hd__a21oi_2 _5403_ (.A1(_3284_),
    .A2(_1332_),
    .B1(_3283_),
    .Y(_1333_));
 sky130_fd_sc_hd__o21bai_1 _5404_ (.A1(_1333_),
    .A2(_1198_),
    .B1_N(_3279_),
    .Y(_1334_));
 sky130_fd_sc_hd__a21oi_2 _5405_ (.A1(_3276_),
    .A2(_1334_),
    .B1(_3275_),
    .Y(_1335_));
 sky130_fd_sc_hd__o21bai_1 _5406_ (.A1(_1331_),
    .A2(_1335_),
    .B1_N(_3271_),
    .Y(_1336_));
 sky130_fd_sc_hd__a21oi_2 _5407_ (.A1(_3268_),
    .A2(_1336_),
    .B1(_3267_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_3432_),
    .B(_3429_),
    .Y(_1338_));
 sky130_fd_sc_hd__a21oi_2 _5409_ (.A1(_3264_),
    .A2(_3431_),
    .B1(_3263_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21ai_2 _5410_ (.A1(_1337_),
    .A2(_1338_),
    .B1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__xor2_4 _5411_ (.A(_3427_),
    .B(net156),
    .X(_3433_));
 sky130_fd_sc_hd__inv_1 _5412_ (.A(_3433_),
    .Y(_3459_));
 sky130_fd_sc_hd__inv_1 _5413_ (.A(_3476_),
    .Y(_1341_));
 sky130_fd_sc_hd__inv_1 _5414_ (.A(_3484_),
    .Y(_1342_));
 sky130_fd_sc_hd__inv_1 _5415_ (.A(_3451_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21o_1 _5416_ (.A1(_2187_),
    .A2(_3457_),
    .B1(_3456_),
    .X(_1344_));
 sky130_fd_sc_hd__a21oi_2 _5417_ (.A1(_1344_),
    .A2(_3455_),
    .B1(_3454_),
    .Y(_1345_));
 sky130_fd_sc_hd__o21bai_1 _5418_ (.A1(_1343_),
    .A2(_1345_),
    .B1_N(_3450_),
    .Y(_1346_));
 sky130_fd_sc_hd__a21oi_2 _5419_ (.A1(_1346_),
    .A2(_3447_),
    .B1(_3446_),
    .Y(_1347_));
 sky130_fd_sc_hd__o21bai_1 _5420_ (.A1(_1342_),
    .A2(_1347_),
    .B1_N(_3483_),
    .Y(_1348_));
 sky130_fd_sc_hd__a21oi_2 _5421_ (.A1(_1348_),
    .A2(_3480_),
    .B1(_3479_),
    .Y(_1349_));
 sky130_fd_sc_hd__o21bai_2 _5422_ (.A1(_1341_),
    .A2(_1349_),
    .B1_N(_3475_),
    .Y(_1350_));
 sky130_fd_sc_hd__a21oi_4 _5423_ (.A1(_3439_),
    .A2(_1350_),
    .B1(_3438_),
    .Y(_1351_));
 sky130_fd_sc_hd__xnor2_4 _5424_ (.A(_3436_),
    .B(net117),
    .Y(_3724_));
 sky130_fd_sc_hd__inv_1 _5425_ (.A(_3724_),
    .Y(_3486_));
 sky130_fd_sc_hd__buf_8 _5426_ (.A(_1316_),
    .X(_3489_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3462_),
    .B(_3489_),
    .Y(_1352_));
 sky130_fd_sc_hd__a21boi_2 _5428_ (.A1(_3517_),
    .A2(_3433_),
    .B1_N(_1352_),
    .Y(_2180_));
 sky130_fd_sc_hd__inv_1 _5429_ (.A(_2180_),
    .Y(_2177_));
 sky130_fd_sc_hd__nor2b_1 _5430_ (.A(_1205_),
    .B_N(_3429_),
    .Y(_1353_));
 sky130_fd_sc_hd__o21a_1 _5431_ (.A1(_3263_),
    .A2(_1353_),
    .B1(_3427_),
    .X(_1354_));
 sky130_fd_sc_hd__nor2_1 _5432_ (.A(_3426_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__xnor2_2 _5433_ (.A(_3468_),
    .B(_1355_),
    .Y(_3469_));
 sky130_fd_sc_hd__xor2_4 _5434_ (.A(_3375_),
    .B(net130),
    .X(_1356_));
 sky130_fd_sc_hd__nor3_1 _5435_ (.A(_3633_),
    .B(_3620_),
    .C(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__nor2b_1 _5436_ (.A(_3641_),
    .B_N(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__nor2b_2 _5437_ (.A(_3649_),
    .B_N(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__nor2b_4 _5438_ (.A(_3657_),
    .B_N(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2b_4 _5439_ (.A_N(_3665_),
    .B(_1360_),
    .Y(_3440_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_1316_),
    .B(_3440_),
    .Y(_1361_));
 sky130_fd_sc_hd__inv_1 _5441_ (.A(_3480_),
    .Y(_1362_));
 sky130_fd_sc_hd__inv_1 _5442_ (.A(_3447_),
    .Y(_1363_));
 sky130_fd_sc_hd__a21o_1 _5443_ (.A1(_2189_),
    .A2(_3455_),
    .B1(_3454_),
    .X(_1364_));
 sky130_fd_sc_hd__a21oi_2 _5444_ (.A1(_3451_),
    .A2(_1364_),
    .B1(_3450_),
    .Y(_1365_));
 sky130_fd_sc_hd__o21bai_1 _5445_ (.A1(_1363_),
    .A2(_1365_),
    .B1_N(_3446_),
    .Y(_1366_));
 sky130_fd_sc_hd__a21oi_2 _5446_ (.A1(_3484_),
    .A2(_1366_),
    .B1(_3483_),
    .Y(_1367_));
 sky130_fd_sc_hd__o21bai_2 _5447_ (.A1(_1362_),
    .A2(_1367_),
    .B1_N(_3479_),
    .Y(_1368_));
 sky130_fd_sc_hd__a21oi_4 _5448_ (.A1(_1368_),
    .A2(net115),
    .B1(_3475_),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2b_4 _5449_ (.A_N(_1369_),
    .B(_3439_),
    .Y(_1370_));
 sky130_fd_sc_hd__nor2_4 _5450_ (.A(_3459_),
    .B(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_1361_),
    .B(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__and2_0 _5452_ (.A(_1316_),
    .B(_3440_),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_4 _5453_ (.A(net179),
    .B(_1370_),
    .Y(_1374_));
 sky130_fd_sc_hd__nand2_1 _5454_ (.A(_1373_),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__a211o_1 _5455_ (.A1(_1372_),
    .A2(_1375_),
    .B1(net124),
    .C1(net148),
    .X(_1376_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_1318_),
    .B(_1374_),
    .Y(_1377_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(net22),
    .B(_1371_),
    .Y(_1378_));
 sky130_fd_sc_hd__a2bb2o_4 _5458_ (.A1_N(net125),
    .A2_N(net135),
    .B1(_1377_),
    .B2(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__a21oi_1 _5459_ (.A1(_3436_),
    .A2(_3438_),
    .B1(_3435_),
    .Y(_1380_));
 sky130_fd_sc_hd__nand3_2 _5460_ (.A(_1376_),
    .B(_1379_),
    .C(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__xor2_2 _5461_ (.A(_3472_),
    .B(_1381_),
    .X(_3728_));
 sky130_fd_sc_hd__xor2_1 _5462_ (.A(_3417_),
    .B(_1300_),
    .X(_1382_));
 sky130_fd_sc_hd__a21o_1 _5463_ (.A1(_3523_),
    .A2(_1382_),
    .B1(_3522_),
    .X(_1383_));
 sky130_fd_sc_hd__a21oi_1 _5464_ (.A1(_3520_),
    .A2(_1383_),
    .B1(_3519_),
    .Y(_1384_));
 sky130_fd_sc_hd__nor2b_1 _5465_ (.A(_1384_),
    .B_N(_3516_),
    .Y(_1385_));
 sky130_fd_sc_hd__o21ai_0 _5466_ (.A1(_3515_),
    .A2(_1385_),
    .B1(_3513_),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2b_1 _5467_ (.A_N(_3512_),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a21oi_1 _5468_ (.A1(_3510_),
    .A2(_1387_),
    .B1(_3509_),
    .Y(_1388_));
 sky130_fd_sc_hd__nor2b_1 _5469_ (.A(_1388_),
    .B_N(_3507_),
    .Y(_1389_));
 sky130_fd_sc_hd__o21ai_0 _5470_ (.A1(_3506_),
    .A2(_1389_),
    .B1(_3504_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2b_1 _5471_ (.A_N(_3503_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a21oi_1 _5472_ (.A1(_3501_),
    .A2(_1391_),
    .B1(_3500_),
    .Y(_1392_));
 sky130_fd_sc_hd__nor2b_1 _5473_ (.A(_1392_),
    .B_N(_3498_),
    .Y(_1393_));
 sky130_fd_sc_hd__o21ai_0 _5474_ (.A1(_3497_),
    .A2(_1393_),
    .B1(_3495_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2b_1 _5475_ (.A_N(_3494_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__a21oi_2 _5476_ (.A1(_3492_),
    .A2(_1395_),
    .B1(_3491_),
    .Y(_1396_));
 sky130_fd_sc_hd__clkbuf_4 _5477_ (.A(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__a21o_2 _5478_ (.A1(_3492_),
    .A2(_1395_),
    .B1(_3491_),
    .X(_1398_));
 sky130_fd_sc_hd__nand2_1 _5479_ (.A(_3488_),
    .B(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__a21boi_2 _5480_ (.A1(net159),
    .A2(_1397_),
    .B1_N(_1399_),
    .Y(_2186_));
 sky130_fd_sc_hd__inv_1 _5481_ (.A(_2186_),
    .Y(_2182_));
 sky130_fd_sc_hd__a21o_1 _5482_ (.A1(_1340_),
    .A2(_3427_),
    .B1(_3426_),
    .X(_1400_));
 sky130_fd_sc_hd__a21oi_2 _5483_ (.A1(_1400_),
    .A2(_3468_),
    .B1(_3467_),
    .Y(_1401_));
 sky130_fd_sc_hd__xnor2_2 _5484_ (.A(_3536_),
    .B(net127),
    .Y(_3537_));
 sky130_fd_sc_hd__nor2_4 _5485_ (.A(_1351_),
    .B(_3459_),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_1402_),
    .B(_1361_),
    .Y(_1403_));
 sky130_fd_sc_hd__nor2_4 _5487_ (.A(net178),
    .B(_1351_),
    .Y(_1404_));
 sky130_fd_sc_hd__nand2_2 _5488_ (.A(_1373_),
    .B(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__a211oi_2 _5489_ (.A1(_1403_),
    .A2(_1405_),
    .B1(net126),
    .C1(net135),
    .Y(_1406_));
 sky130_fd_sc_hd__nand2_1 _5490_ (.A(_1318_),
    .B(_1404_),
    .Y(_1407_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(net22),
    .B(_1402_),
    .Y(_1408_));
 sky130_fd_sc_hd__a2bb2oi_1 _5492_ (.A1_N(net125),
    .A2_N(net135),
    .B1(_1407_),
    .B2(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2b_1 _5493_ (.A_N(_3435_),
    .B(_3540_),
    .Y(_1410_));
 sky130_fd_sc_hd__or4_4 _5494_ (.A(_3471_),
    .B(_1406_),
    .C(_1409_),
    .D(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__nor2b_1 _5495_ (.A(_3540_),
    .B_N(_3472_),
    .Y(_1412_));
 sky130_fd_sc_hd__o21ai_1 _5496_ (.A1(_1409_),
    .A2(_1406_),
    .B1(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__inv_1 _5497_ (.A(_3540_),
    .Y(_1414_));
 sky130_fd_sc_hd__nor3_1 _5498_ (.A(_3472_),
    .B(_1414_),
    .C(_3471_),
    .Y(_1415_));
 sky130_fd_sc_hd__a221oi_2 _5499_ (.A1(_1414_),
    .A2(_3471_),
    .B1(_1412_),
    .B2(_3435_),
    .C1(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand3_2 _5500_ (.A(_1413_),
    .B(_1411_),
    .C(_1416_),
    .Y(_3732_));
 sky130_fd_sc_hd__o21ai_0 _5501_ (.A1(_3426_),
    .A2(_1354_),
    .B1(_3468_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2b_1 _5502_ (.A_N(_3467_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__a21oi_2 _5503_ (.A1(_3536_),
    .A2(_1418_),
    .B1(_3535_),
    .Y(_1419_));
 sky130_fd_sc_hd__xnor2_2 _5504_ (.A(_3552_),
    .B(_1419_),
    .Y(_3554_));
 sky130_fd_sc_hd__nor3b_1 _5505_ (.A(_3471_),
    .B(_3539_),
    .C_N(_1380_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand3_1 _5506_ (.A(net175),
    .B(_1379_),
    .C(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nor2_1 _5507_ (.A(_3472_),
    .B(_3471_),
    .Y(_1422_));
 sky130_fd_sc_hd__o21bai_1 _5508_ (.A1(_1414_),
    .A2(_1422_),
    .B1_N(_3539_),
    .Y(_1423_));
 sky130_fd_sc_hd__nand2_2 _5509_ (.A(_1421_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__xnor2_4 _5510_ (.A(_3556_),
    .B(_1424_),
    .Y(_3736_));
 sky130_fd_sc_hd__nor2b_1 _5511_ (.A(_1401_),
    .B_N(_3536_),
    .Y(_1425_));
 sky130_fd_sc_hd__o21ai_1 _5512_ (.A1(_3535_),
    .A2(_1425_),
    .B1(_3552_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2b_2 _5513_ (.A_N(_3551_),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__xor2_4 _5514_ (.A(_3568_),
    .B(net141),
    .X(_3569_));
 sky130_fd_sc_hd__xnor3_1 _5515_ (.A(_3198_),
    .B(_1324_),
    .C(net136),
    .X(_1428_));
 sky130_fd_sc_hd__a21o_1 _5516_ (.A1(_1320_),
    .A2(_1321_),
    .B1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__nand3_2 _5517_ (.A(_1320_),
    .B(_1321_),
    .C(_1428_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand3_4 _5518_ (.A(net211),
    .B(_1429_),
    .C(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__or3_1 _5519_ (.A(net123),
    .B(net148),
    .C(_1361_),
    .X(_1432_));
 sky130_fd_sc_hd__buf_4 _5520_ (.A(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__and3_1 _5521_ (.A(_3472_),
    .B(_3540_),
    .C(_1402_),
    .X(_1434_));
 sky130_fd_sc_hd__nand3_1 _5522_ (.A(_1431_),
    .B(_1433_),
    .C(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand3_1 _5523_ (.A(_3472_),
    .B(_3540_),
    .C(_1404_),
    .Y(_1436_));
 sky130_fd_sc_hd__a21o_1 _5524_ (.A1(_1431_),
    .A2(_1433_),
    .B1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__a21o_1 _5525_ (.A1(_3472_),
    .A2(_3435_),
    .B1(_3471_),
    .X(_1438_));
 sky130_fd_sc_hd__a21oi_1 _5526_ (.A1(_3540_),
    .A2(_1438_),
    .B1(_3539_),
    .Y(_1439_));
 sky130_fd_sc_hd__inv_1 _5527_ (.A(_3556_),
    .Y(_1440_));
 sky130_fd_sc_hd__a31oi_1 _5528_ (.A1(_1435_),
    .A2(_1437_),
    .A3(_1439_),
    .B1(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__or2_0 _5529_ (.A(_3572_),
    .B(_3555_),
    .X(_1442_));
 sky130_fd_sc_hd__a21o_1 _5530_ (.A1(_3540_),
    .A2(_1438_),
    .B1(_3539_),
    .X(_1443_));
 sky130_fd_sc_hd__nor2_1 _5531_ (.A(_3555_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__or2_0 _5532_ (.A(_3556_),
    .B(_3555_),
    .X(_1445_));
 sky130_fd_sc_hd__nand2_1 _5533_ (.A(_3572_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__a31oi_2 _5534_ (.A1(_1435_),
    .A2(_1437_),
    .A3(_1444_),
    .B1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__o21ba_1 _5535_ (.A1(_1441_),
    .A2(_1442_),
    .B1_N(_1447_),
    .X(_3740_));
 sky130_fd_sc_hd__inv_1 _5536_ (.A(_3552_),
    .Y(_1448_));
 sky130_fd_sc_hd__o21bai_1 _5537_ (.A1(_1448_),
    .A2(_1419_),
    .B1_N(_3551_),
    .Y(_1449_));
 sky130_fd_sc_hd__a21oi_2 _5538_ (.A1(_3568_),
    .A2(_1449_),
    .B1(_3567_),
    .Y(_1450_));
 sky130_fd_sc_hd__xnor2_4 _5539_ (.A(_3584_),
    .B(_1450_),
    .Y(_3585_));
 sky130_fd_sc_hd__nand2_1 _5540_ (.A(_3556_),
    .B(_3572_),
    .Y(_1451_));
 sky130_fd_sc_hd__inv_1 _5541_ (.A(_3588_),
    .Y(_1452_));
 sky130_fd_sc_hd__a2111o_1 _5542_ (.A1(_1423_),
    .A2(_1421_),
    .B1(_1452_),
    .C1(_3555_),
    .D1(_3571_),
    .X(_1453_));
 sky130_fd_sc_hd__or4_1 _5543_ (.A(_3556_),
    .B(_1452_),
    .C(_3555_),
    .D(_3571_),
    .X(_1454_));
 sky130_fd_sc_hd__nor2b_1 _5544_ (.A(_3588_),
    .B_N(_3571_),
    .Y(_1455_));
 sky130_fd_sc_hd__a31oi_1 _5545_ (.A1(_3572_),
    .A2(_1452_),
    .A3(_3555_),
    .B1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__o311a_1 _5546_ (.A1(_3572_),
    .A2(_1452_),
    .A3(_3571_),
    .B1(_1454_),
    .C1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__o311ai_4 _5547_ (.A1(_3588_),
    .A2(_1424_),
    .A3(_1451_),
    .B1(_1453_),
    .C1(_1457_),
    .Y(_3743_));
 sky130_fd_sc_hd__nor3_1 _5548_ (.A(_3372_),
    .B(_3328_),
    .C(_3376_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand2b_1 _5549_ (.A_N(_3324_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__or2_0 _5550_ (.A(_3365_),
    .B(_3368_),
    .X(_1460_));
 sky130_fd_sc_hd__or3_1 _5551_ (.A(_3361_),
    .B(_1459_),
    .C(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__or3_4 _5552_ (.A(net139),
    .B(_1128_),
    .C(_1324_),
    .X(_1462_));
 sky130_fd_sc_hd__o21ai_2 _5553_ (.A1(net139),
    .A2(_1128_),
    .B1(_1324_),
    .Y(_1463_));
 sky130_fd_sc_hd__o2111ai_4 _5554_ (.A1(_3321_),
    .A2(_1461_),
    .B1(_1462_),
    .C1(_1463_),
    .D1(_1185_),
    .Y(_1464_));
 sky130_fd_sc_hd__a21o_2 _5555_ (.A1(_1463_),
    .A2(_1462_),
    .B1(_1185_),
    .X(_1465_));
 sky130_fd_sc_hd__or2_2 _5556_ (.A(_1233_),
    .B(_1240_),
    .X(_3311_));
 sky130_fd_sc_hd__a21o_1 _5557_ (.A1(_3568_),
    .A2(_1427_),
    .B1(_3567_),
    .X(_1466_));
 sky130_fd_sc_hd__a21oi_2 _5558_ (.A1(_3584_),
    .A2(_1466_),
    .B1(_3583_),
    .Y(_1467_));
 sky130_fd_sc_hd__xor3_2 _5559_ (.A(_3311_),
    .B(_1467_),
    .C(_1244_),
    .X(_1468_));
 sky130_fd_sc_hd__a21oi_4 _5560_ (.A1(_1464_),
    .A2(_1465_),
    .B1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__and3_4 _5561_ (.A(_1464_),
    .B(_1465_),
    .C(_1468_),
    .X(_1470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__nor2_8 _5563_ (.A(_1469_),
    .B(_1470_),
    .Y(_1472_));
 sky130_fd_sc_hd__clkinv_4 _5564_ (.A(_1472_),
    .Y(_3606_));
 sky130_fd_sc_hd__nor3b_1 _5565_ (.A(_3469_),
    .B(_3537_),
    .C_N(_3461_),
    .Y(_1473_));
 sky130_fd_sc_hd__nor3b_1 _5566_ (.A(_3554_),
    .B(_3569_),
    .C_N(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nor2_1 _5567_ (.A(net21),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__o21ai_0 _5568_ (.A1(_3585_),
    .A2(_1475_),
    .B1(_3489_),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_4 _5569_ (.A(net188),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a21oi_1 _5570_ (.A1(net27),
    .A2(_1472_),
    .B1(_1477_),
    .Y(_3621_));
 sky130_fd_sc_hd__and2_0 _5571_ (.A(_3442_),
    .B(_3489_),
    .X(_1478_));
 sky130_fd_sc_hd__a31oi_4 _5572_ (.A1(net21),
    .A2(_1429_),
    .A3(_1430_),
    .B1(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__xnor2_4 _5573_ (.A(net29),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nor3_1 _5574_ (.A(_3555_),
    .B(_3571_),
    .C(_1443_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand3_1 _5575_ (.A(_1435_),
    .B(_1437_),
    .C(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__a21oi_1 _5576_ (.A1(_3572_),
    .A2(_1445_),
    .B1(_3571_),
    .Y(_1483_));
 sky130_fd_sc_hd__inv_1 _5577_ (.A(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand4_2 _5578_ (.A(_3588_),
    .B(_1480_),
    .C(_1482_),
    .D(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__or4_2 _5579_ (.A(_3571_),
    .B(_3587_),
    .C(_1447_),
    .D(_1480_),
    .X(_1486_));
 sky130_fd_sc_hd__nor3_1 _5580_ (.A(_3588_),
    .B(_3587_),
    .C(_1480_),
    .Y(_1487_));
 sky130_fd_sc_hd__a21oi_2 _5581_ (.A1(_3587_),
    .A2(_1480_),
    .B1(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand3_1 _5582_ (.A(_1485_),
    .B(_1486_),
    .C(_1488_),
    .Y(_3598_));
 sky130_fd_sc_hd__or3_1 _5583_ (.A(_3292_),
    .B(_3433_),
    .C(_3469_),
    .X(_1489_));
 sky130_fd_sc_hd__or3_4 _5584_ (.A(_3537_),
    .B(_3554_),
    .C(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__nor3_4 _5585_ (.A(_3569_),
    .B(_1490_),
    .C(_3585_),
    .Y(_1491_));
 sky130_fd_sc_hd__nor2_1 _5586_ (.A(net21),
    .B(net195),
    .Y(_1492_));
 sky130_fd_sc_hd__mux2i_4 _5587_ (.A0(net21),
    .A1(_1492_),
    .S(net192),
    .Y(_3640_));
 sky130_fd_sc_hd__nor2b_1 _5588_ (.A(_2176_),
    .B_N(_3464_),
    .Y(_1493_));
 sky130_fd_sc_hd__o21ai_1 _5589_ (.A1(_3463_),
    .A2(_1493_),
    .B1(_3532_),
    .Y(_1494_));
 sky130_fd_sc_hd__nand2b_1 _5590_ (.A_N(_3531_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__a21o_1 _5591_ (.A1(_1495_),
    .A2(_3548_),
    .B1(_3547_),
    .X(_1496_));
 sky130_fd_sc_hd__a21o_1 _5592_ (.A1(_1496_),
    .A2(_3564_),
    .B1(_3563_),
    .X(_1497_));
 sky130_fd_sc_hd__a21o_1 _5593_ (.A1(_1497_),
    .A2(_3580_),
    .B1(_3579_),
    .X(_1498_));
 sky130_fd_sc_hd__a21o_1 _5594_ (.A1(_1498_),
    .A2(_3596_),
    .B1(_3595_),
    .X(_1499_));
 sky130_fd_sc_hd__a21o_1 _5595_ (.A1(_3612_),
    .A2(_1499_),
    .B1(_3611_),
    .X(_1500_));
 sky130_fd_sc_hd__a21o_1 _5596_ (.A1(_1500_),
    .A2(_3623_),
    .B1(_3622_),
    .X(_1501_));
 sky130_fd_sc_hd__xnor2_4 _5597_ (.A(net145),
    .B(_1356_),
    .Y(_1502_));
 sky130_fd_sc_hd__xnor2_4 _5598_ (.A(_3640_),
    .B(_1502_),
    .Y(_3629_));
 sky130_fd_sc_hd__inv_1 _5599_ (.A(_3629_),
    .Y(_3673_));
 sky130_fd_sc_hd__or3_4 _5600_ (.A(_3724_),
    .B(_3732_),
    .C(net157),
    .X(_1503_));
 sky130_fd_sc_hd__or4_4 _5601_ (.A(_3736_),
    .B(_3740_),
    .C(_1503_),
    .D(_3743_),
    .X(_1504_));
 sky130_fd_sc_hd__a31oi_4 _5602_ (.A1(_1485_),
    .A2(_1486_),
    .A3(_1488_),
    .B1(_1397_),
    .Y(_1505_));
 sky130_fd_sc_hd__and4_1 _5603_ (.A(_1396_),
    .B(_1485_),
    .C(_1486_),
    .D(_1488_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_2 _5604_ (.A(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__a21oi_1 _5605_ (.A1(net180),
    .A2(_1505_),
    .B1(_1507_),
    .Y(_3628_));
 sky130_fd_sc_hd__a21oi_1 _5606_ (.A1(net27),
    .A2(_1472_),
    .B1(_1477_),
    .Y(_3632_));
 sky130_fd_sc_hd__nor2b_1 _5607_ (.A(_2178_),
    .B_N(_3532_),
    .Y(_1508_));
 sky130_fd_sc_hd__o21ai_1 _5608_ (.A1(_1508_),
    .A2(_3531_),
    .B1(_3548_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2b_1 _5609_ (.A_N(_3547_),
    .B(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__a21o_1 _5610_ (.A1(_1510_),
    .A2(_3564_),
    .B1(_3563_),
    .X(_1511_));
 sky130_fd_sc_hd__a21o_1 _5611_ (.A1(_1511_),
    .A2(_3580_),
    .B1(_3579_),
    .X(_1512_));
 sky130_fd_sc_hd__a21o_1 _5612_ (.A1(_1512_),
    .A2(_3596_),
    .B1(_3595_),
    .X(_1513_));
 sky130_fd_sc_hd__a21o_1 _5613_ (.A1(_3612_),
    .A2(_1513_),
    .B1(_3611_),
    .X(_1514_));
 sky130_fd_sc_hd__a21o_1 _5614_ (.A1(_1514_),
    .A2(_3623_),
    .B1(_3622_),
    .X(_1515_));
 sky130_fd_sc_hd__or2_1 _5615_ (.A(_1316_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__nor3_4 _5616_ (.A(net149),
    .B(net195),
    .C(_1515_),
    .Y(_1517_));
 sky130_fd_sc_hd__o21ai_2 _5617_ (.A1(net203),
    .A2(net199),
    .B1(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_0 _5618_ (.A(_1356_),
    .B(_1515_),
    .X(_1519_));
 sky130_fd_sc_hd__o211a_1 _5619_ (.A1(net193),
    .A2(_1516_),
    .B1(_1518_),
    .C1(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__nor3_1 _5620_ (.A(net212),
    .B(_1356_),
    .C(_1491_),
    .Y(_1521_));
 sky130_fd_sc_hd__nor2_1 _5621_ (.A(net22),
    .B(_1356_),
    .Y(_1522_));
 sky130_fd_sc_hd__mux2i_1 _5622_ (.A0(_1521_),
    .A1(_1522_),
    .S(net29),
    .Y(_1523_));
 sky130_fd_sc_hd__inv_1 _5623_ (.A(_3635_),
    .Y(_1524_));
 sky130_fd_sc_hd__a21oi_2 _5624_ (.A1(_1523_),
    .A2(_1520_),
    .B1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand3_2 _5625_ (.A(net272),
    .B(_1524_),
    .C(_1523_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2b_4 _5626_ (.A_N(_1525_),
    .B(_1526_),
    .Y(_3636_));
 sky130_fd_sc_hd__nand4_2 _5627_ (.A(_3487_),
    .B(_1411_),
    .C(net122),
    .D(_1416_),
    .Y(_1527_));
 sky130_fd_sc_hd__or4_4 _5628_ (.A(_3736_),
    .B(_1527_),
    .C(_3743_),
    .D(_3740_),
    .X(_3597_));
 sky130_fd_sc_hd__a21oi_1 _5629_ (.A1(_1505_),
    .A2(_3597_),
    .B1(_1507_),
    .Y(_3637_));
 sky130_fd_sc_hd__inv_1 _5630_ (.A(_1491_),
    .Y(_3605_));
 sky130_fd_sc_hd__nand2_2 _5631_ (.A(_1356_),
    .B(_1501_),
    .Y(_1528_));
 sky130_fd_sc_hd__o2111a_2 _5632_ (.A1(net204),
    .A2(net205),
    .B1(_3605_),
    .C1(net22),
    .D1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__nand2_2 _5633_ (.A(net147),
    .B(net206),
    .Y(_1530_));
 sky130_fd_sc_hd__nor3_4 _5634_ (.A(net189),
    .B(_1530_),
    .C(net121),
    .Y(_1531_));
 sky130_fd_sc_hd__o21ai_2 _5635_ (.A1(net145),
    .A2(_1356_),
    .B1(_3635_),
    .Y(_1532_));
 sky130_fd_sc_hd__inv_1 _5636_ (.A(_3634_),
    .Y(_1533_));
 sky130_fd_sc_hd__o31ai_4 _5637_ (.A1(_1529_),
    .A2(net143),
    .A3(net146),
    .B1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__xnor2_4 _5638_ (.A(_3643_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__inv_1 _5639_ (.A(_1535_),
    .Y(_3645_));
 sky130_fd_sc_hd__a21oi_1 _5640_ (.A1(net181),
    .A2(_1505_),
    .B1(_1507_),
    .Y(_3644_));
 sky130_fd_sc_hd__a21oi_1 _5641_ (.A1(net27),
    .A2(net29),
    .B1(_1477_),
    .Y(_3648_));
 sky130_fd_sc_hd__o211ai_2 _5642_ (.A1(net193),
    .A2(net237),
    .B1(_1519_),
    .C1(_1518_),
    .Y(_1536_));
 sky130_fd_sc_hd__mux2_1 _5643_ (.A0(_1521_),
    .A1(_1522_),
    .S(net29),
    .X(_1537_));
 sky130_fd_sc_hd__nand2_1 _5644_ (.A(_3635_),
    .B(_3643_),
    .Y(_1538_));
 sky130_fd_sc_hd__a21oi_1 _5645_ (.A1(_3643_),
    .A2(_3634_),
    .B1(_3642_),
    .Y(_1539_));
 sky130_fd_sc_hd__o31a_4 _5646_ (.A1(_1538_),
    .A2(_1537_),
    .A3(_1536_),
    .B1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__xnor2_4 _5647_ (.A(_3651_),
    .B(_1540_),
    .Y(_3653_));
 sky130_fd_sc_hd__a21oi_1 _5648_ (.A1(_1505_),
    .A2(_3597_),
    .B1(_1507_),
    .Y(_3652_));
 sky130_fd_sc_hd__mux2i_1 _5649_ (.A0(net27),
    .A1(_1492_),
    .S(_3606_),
    .Y(_3656_));
 sky130_fd_sc_hd__nor3_2 _5650_ (.A(net223),
    .B(_1531_),
    .C(_1532_),
    .Y(_1541_));
 sky130_fd_sc_hd__nor3_1 _5651_ (.A(_3643_),
    .B(_3642_),
    .C(_3650_),
    .Y(_1542_));
 sky130_fd_sc_hd__nor2_1 _5652_ (.A(_3651_),
    .B(_3650_),
    .Y(_1543_));
 sky130_fd_sc_hd__nor2_1 _5653_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__o41ai_4 _5654_ (.A1(_3634_),
    .A2(_1541_),
    .A3(_3650_),
    .A4(_3642_),
    .B1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__xnor2_4 _5655_ (.A(_3659_),
    .B(net110),
    .Y(_3661_));
 sky130_fd_sc_hd__a21oi_1 _5656_ (.A1(net180),
    .A2(_1505_),
    .B1(_1507_),
    .Y(_3660_));
 sky130_fd_sc_hd__a21oi_1 _5657_ (.A1(net27),
    .A2(net188),
    .B1(_1477_),
    .Y(_3664_));
 sky130_fd_sc_hd__nand2_1 _5658_ (.A(_3651_),
    .B(_3659_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor3b_1 _5659_ (.A(_3650_),
    .B(_3658_),
    .C_N(_3667_),
    .Y(_1547_));
 sky130_fd_sc_hd__o311ai_4 _5660_ (.A1(_1536_),
    .A2(_1537_),
    .A3(_1538_),
    .B1(_1539_),
    .C1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__nor4b_1 _5661_ (.A(_3651_),
    .B(_3650_),
    .C(_3658_),
    .D_N(_3667_),
    .Y(_1549_));
 sky130_fd_sc_hd__nor3b_1 _5662_ (.A(_3659_),
    .B(_3658_),
    .C_N(_3667_),
    .Y(_1550_));
 sky130_fd_sc_hd__inv_1 _5663_ (.A(_3658_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand3b_1 _5664_ (.A_N(_3667_),
    .B(_3650_),
    .C(_3659_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21ai_0 _5665_ (.A1(_3667_),
    .A2(_1551_),
    .B1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__nor3_1 _5666_ (.A(_1549_),
    .B(_1550_),
    .C(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__o311ai_4 _5667_ (.A1(_3667_),
    .A2(_1540_),
    .A3(_1546_),
    .B1(_1548_),
    .C1(_1554_),
    .Y(_3669_));
 sky130_fd_sc_hd__buf_2 _5668_ (.A(_1398_),
    .X(_1555_));
 sky130_fd_sc_hd__a21oi_1 _5669_ (.A1(_3599_),
    .A2(_1555_),
    .B1(_1507_),
    .Y(_3668_));
 sky130_fd_sc_hd__o21ai_1 _5670_ (.A1(_1469_),
    .A2(_1470_),
    .B1(net21),
    .Y(_1556_));
 sky130_fd_sc_hd__nand2b_1 _5671_ (.A_N(_3607_),
    .B(_3489_),
    .Y(_1557_));
 sky130_fd_sc_hd__nand3_1 _5672_ (.A(_1330_),
    .B(_1556_),
    .C(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__a21o_1 _5673_ (.A1(_1556_),
    .A2(_1557_),
    .B1(_1330_),
    .X(_1559_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_1558_),
    .B(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_3659_),
    .B(_3667_),
    .Y(_1561_));
 sky130_fd_sc_hd__and2_0 _5676_ (.A(_3667_),
    .B(_3658_),
    .X(_1562_));
 sky130_fd_sc_hd__o211ai_1 _5677_ (.A1(_3666_),
    .A2(_1562_),
    .B1(_1559_),
    .C1(_1558_),
    .Y(_1563_));
 sky130_fd_sc_hd__o31a_1 _5678_ (.A1(_1561_),
    .A2(_1560_),
    .A3(net111),
    .B1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__nor2_1 _5679_ (.A(_3658_),
    .B(_3666_),
    .Y(_1565_));
 sky130_fd_sc_hd__or2_0 _5680_ (.A(_3659_),
    .B(_3658_),
    .X(_1566_));
 sky130_fd_sc_hd__a221oi_2 _5681_ (.A1(_1558_),
    .A2(_1559_),
    .B1(_1566_),
    .B2(_3667_),
    .C1(_3666_),
    .Y(_1567_));
 sky130_fd_sc_hd__a31oi_4 _5682_ (.A1(net112),
    .A2(_1560_),
    .A3(_1565_),
    .B1(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__and2_2 _5683_ (.A(_1564_),
    .B(_1568_),
    .X(_3705_));
 sky130_fd_sc_hd__clkinv_4 _5684_ (.A(_3636_),
    .Y(_3672_));
 sky130_fd_sc_hd__inv_4 _5685_ (.A(net239),
    .Y(_3679_));
 sky130_fd_sc_hd__inv_1 _5686_ (.A(net78),
    .Y(_3680_));
 sky130_fd_sc_hd__inv_1 _5687_ (.A(_2331_),
    .Y(_2094_));
 sky130_fd_sc_hd__inv_1 _5688_ (.A(_2199_),
    .Y(_2083_));
 sky130_fd_sc_hd__inv_1 _5689_ (.A(_2103_),
    .Y(_2118_));
 sky130_fd_sc_hd__inv_1 _5690_ (.A(_2135_),
    .Y(_2142_));
 sky130_fd_sc_hd__inv_1 _5691_ (.A(_2173_),
    .Y(_2175_));
 sky130_fd_sc_hd__inv_1 _5692_ (.A(net30),
    .Y(_2195_));
 sky130_fd_sc_hd__inv_1 _5693_ (.A(net37),
    .Y(_2078_));
 sky130_fd_sc_hd__inv_1 _5694_ (.A(net39),
    .Y(_2209_));
 sky130_fd_sc_hd__inv_1 _5695_ (.A(net38),
    .Y(_2217_));
 sky130_fd_sc_hd__or2_0 _5696_ (.A(_3685_),
    .B(_0004_),
    .X(_1569_));
 sky130_fd_sc_hd__nand2b_4 _5697_ (.A_N(net70),
    .B(_2472_),
    .Y(_1570_));
 sky130_fd_sc_hd__or4_4 _5698_ (.A(net73),
    .B(net72),
    .C(_1570_),
    .D(net71),
    .X(_1571_));
 sky130_fd_sc_hd__o31ai_4 _5699_ (.A1(net74),
    .A2(_1571_),
    .A3(_0005_),
    .B1(_0040_),
    .Y(_1572_));
 sky130_fd_sc_hd__o21ai_2 _5700_ (.A1(_0003_),
    .A2(_1569_),
    .B1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__xnor2_2 _5701_ (.A(_1573_),
    .B(_3683_),
    .Y(_2090_));
 sky130_fd_sc_hd__inv_1 _5702_ (.A(net41),
    .Y(_2239_));
 sky130_fd_sc_hd__inv_1 _5703_ (.A(net40),
    .Y(_2247_));
 sky130_fd_sc_hd__inv_1 _5704_ (.A(net42),
    .Y(_2255_));
 sky130_fd_sc_hd__o21ai_0 _5705_ (.A1(net64),
    .A2(net63),
    .B1(_0041_),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_1 _5706_ (.A(_1572_),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__xor2_1 _5707_ (.A(net65),
    .B(_1575_),
    .X(_2287_));
 sky130_fd_sc_hd__o21ai_0 _5708_ (.A1(net63),
    .A2(_0039_),
    .B1(_0041_),
    .Y(_1576_));
 sky130_fd_sc_hd__xnor2_1 _5709_ (.A(net64),
    .B(_1576_),
    .Y(_2290_));
 sky130_fd_sc_hd__xnor2_1 _5710_ (.A(net63),
    .B(_1572_),
    .Y(_2293_));
 sky130_fd_sc_hd__o31ai_1 _5711_ (.A1(net76),
    .A2(net75),
    .A3(_0038_),
    .B1(_0041_),
    .Y(_1577_));
 sky130_fd_sc_hd__xnor2_1 _5712_ (.A(net77),
    .B(_1577_),
    .Y(_2296_));
 sky130_fd_sc_hd__o31ai_1 _5713_ (.A1(net75),
    .A2(net74),
    .A3(_1571_),
    .B1(_0041_),
    .Y(_1578_));
 sky130_fd_sc_hd__xnor2_1 _5714_ (.A(net76),
    .B(_1578_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _5715_ (.A(_0038_),
    .B(_0041_),
    .Y(_1579_));
 sky130_fd_sc_hd__xnor2_1 _5716_ (.A(net75),
    .B(_1579_),
    .Y(_2302_));
 sky130_fd_sc_hd__nand2_1 _5717_ (.A(_0041_),
    .B(_1571_),
    .Y(_1580_));
 sky130_fd_sc_hd__xnor2_1 _5718_ (.A(net74),
    .B(_1580_),
    .Y(_2305_));
 sky130_fd_sc_hd__nor2_1 _5719_ (.A(net72),
    .B(net71),
    .Y(_1581_));
 sky130_fd_sc_hd__a21oi_1 _5720_ (.A1(_0000_),
    .A2(_1581_),
    .B1(_1569_),
    .Y(_1582_));
 sky130_fd_sc_hd__xor2_1 _5721_ (.A(net73),
    .B(_1582_),
    .X(_2308_));
 sky130_fd_sc_hd__o21ai_0 _5722_ (.A1(net71),
    .A2(_1570_),
    .B1(_0041_),
    .Y(_1583_));
 sky130_fd_sc_hd__xnor2_1 _5723_ (.A(net72),
    .B(_1583_),
    .Y(_2311_));
 sky130_fd_sc_hd__nor2_1 _5724_ (.A(_0000_),
    .B(_1569_),
    .Y(_1584_));
 sky130_fd_sc_hd__xor2_2 _5725_ (.A(net71),
    .B(_1584_),
    .X(_2107_));
 sky130_fd_sc_hd__nor2_1 _5726_ (.A(_2088_),
    .B(_2091_),
    .Y(_1585_));
 sky130_fd_sc_hd__nand2_1 _5727_ (.A(_2087_),
    .B(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__o31ai_1 _5728_ (.A1(_2085_),
    .A2(_0033_),
    .A3(_0015_),
    .B1(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__nand3b_1 _5729_ (.A_N(_2085_),
    .B(_0033_),
    .C(_2091_),
    .Y(_1588_));
 sky130_fd_sc_hd__o311ai_0 _5730_ (.A1(_2088_),
    .A2(_2087_),
    .A3(_2091_),
    .B1(_1588_),
    .C1(_0032_),
    .Y(_1589_));
 sky130_fd_sc_hd__o21ai_0 _5731_ (.A1(_0032_),
    .A2(_1587_),
    .B1(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__o21ai_0 _5732_ (.A1(_2272_),
    .A2(_1590_),
    .B1(_0125_),
    .Y(_1591_));
 sky130_fd_sc_hd__xnor2_1 _5733_ (.A(_2268_),
    .B(_1591_),
    .Y(_2316_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(_2329_),
    .B(net15),
    .Y(_1592_));
 sky130_fd_sc_hd__xor2_1 _5735_ (.A(_2416_),
    .B(_1592_),
    .X(_2324_));
 sky130_fd_sc_hd__inv_1 _5736_ (.A(net43),
    .Y(_2339_));
 sky130_fd_sc_hd__inv_1 _5737_ (.A(net44),
    .Y(_2347_));
 sky130_fd_sc_hd__inv_1 _5738_ (.A(net31),
    .Y(_2363_));
 sky130_fd_sc_hd__inv_1 _5739_ (.A(net45),
    .Y(_2371_));
 sky130_fd_sc_hd__or2_0 _5740_ (.A(_0025_),
    .B(_0113_),
    .X(_1593_));
 sky130_fd_sc_hd__nand3_1 _5741_ (.A(net172),
    .B(_0029_),
    .C(_0090_),
    .Y(_1594_));
 sky130_fd_sc_hd__o21ai_2 _5742_ (.A1(_0010_),
    .A2(_1593_),
    .B1(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_2 _5743_ (.A(_2232_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__o21ai_0 _5744_ (.A1(_0682_),
    .A2(_1596_),
    .B1(_0125_),
    .Y(_1597_));
 sky130_fd_sc_hd__xnor2_1 _5745_ (.A(_2502_),
    .B(_1597_),
    .Y(_2383_));
 sky130_fd_sc_hd__nor2_1 _5746_ (.A(_0680_),
    .B(_0681_),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_0 _5747_ (.A1(_1598_),
    .A2(_0688_),
    .B1(_0125_),
    .Y(_1599_));
 sky130_fd_sc_hd__xnor2_1 _5748_ (.A(_2506_),
    .B(_1599_),
    .Y(_2387_));
 sky130_fd_sc_hd__nor3_1 _5749_ (.A(_0015_),
    .B(_0064_),
    .C(_0078_),
    .Y(_1600_));
 sky130_fd_sc_hd__a31oi_1 _5750_ (.A1(_0016_),
    .A2(_0053_),
    .A3(_0214_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__o21ai_0 _5751_ (.A1(_1596_),
    .A2(_1601_),
    .B1(_0125_),
    .Y(_1602_));
 sky130_fd_sc_hd__xnor2_1 _5752_ (.A(_2356_),
    .B(_1602_),
    .Y(_2391_));
 sky130_fd_sc_hd__o21ai_0 _5753_ (.A1(_2264_),
    .A2(_0688_),
    .B1(_0125_),
    .Y(_1603_));
 sky130_fd_sc_hd__xnor2_1 _5754_ (.A(_2360_),
    .B(_1603_),
    .Y(_2395_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_0115_),
    .B(_1596_),
    .Y(_1604_));
 sky130_fd_sc_hd__xnor2_1 _5756_ (.A(_2264_),
    .B(_1604_),
    .Y(_2399_));
 sky130_fd_sc_hd__inv_1 _5757_ (.A(_2289_),
    .Y(_1605_));
 sky130_fd_sc_hd__inv_1 _5758_ (.A(_2295_),
    .Y(_1606_));
 sky130_fd_sc_hd__a21o_1 _5759_ (.A1(_2108_),
    .A2(_2313_),
    .B1(_2312_),
    .X(_1607_));
 sky130_fd_sc_hd__a21oi_1 _5760_ (.A1(_2310_),
    .A2(_1607_),
    .B1(_2309_),
    .Y(_1608_));
 sky130_fd_sc_hd__o21bai_1 _5761_ (.A1(_0145_),
    .A2(_1608_),
    .B1_N(_2306_),
    .Y(_1609_));
 sky130_fd_sc_hd__a21oi_1 _5762_ (.A1(_2304_),
    .A2(_1609_),
    .B1(_2303_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21bai_1 _5763_ (.A1(_0146_),
    .A2(_1610_),
    .B1_N(_2300_),
    .Y(_1611_));
 sky130_fd_sc_hd__a21oi_1 _5764_ (.A1(_2298_),
    .A2(_1611_),
    .B1(_2297_),
    .Y(_1612_));
 sky130_fd_sc_hd__o21ai_0 _5765_ (.A1(_1606_),
    .A2(_1612_),
    .B1(_0141_),
    .Y(_1613_));
 sky130_fd_sc_hd__a21oi_1 _5766_ (.A1(_2292_),
    .A2(_1613_),
    .B1(_2291_),
    .Y(_1614_));
 sky130_fd_sc_hd__o21bai_1 _5767_ (.A1(_1605_),
    .A2(_1614_),
    .B1_N(_2288_),
    .Y(_1615_));
 sky130_fd_sc_hd__a21oi_1 _5768_ (.A1(_2286_),
    .A2(_1615_),
    .B1(_2285_),
    .Y(_1616_));
 sky130_fd_sc_hd__xor2_1 _5769_ (.A(_0155_),
    .B(_1616_),
    .X(_2433_));
 sky130_fd_sc_hd__nor2_1 _5770_ (.A(_2291_),
    .B(_0154_),
    .Y(_1617_));
 sky130_fd_sc_hd__nor2_1 _5771_ (.A(_1605_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nor2_1 _5772_ (.A(_2288_),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__xnor2_1 _5773_ (.A(_2286_),
    .B(_1619_),
    .Y(_2436_));
 sky130_fd_sc_hd__xnor2_1 _5774_ (.A(_2289_),
    .B(_1614_),
    .Y(_2439_));
 sky130_fd_sc_hd__a21oi_1 _5775_ (.A1(_0149_),
    .A2(_0152_),
    .B1(_1606_),
    .Y(_1620_));
 sky130_fd_sc_hd__nor3_1 _5776_ (.A(_2292_),
    .B(_2294_),
    .C(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__nor2_1 _5777_ (.A(_0154_),
    .B(_1621_),
    .Y(_2442_));
 sky130_fd_sc_hd__xnor2_1 _5778_ (.A(_2295_),
    .B(_1612_),
    .Y(_2446_));
 sky130_fd_sc_hd__nor2_1 _5779_ (.A(_2309_),
    .B(_0144_),
    .Y(_1622_));
 sky130_fd_sc_hd__nor2_1 _5780_ (.A(_0145_),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a31oi_1 _5781_ (.A1(_2304_),
    .A2(_2301_),
    .A3(_1623_),
    .B1(_0151_),
    .Y(_1624_));
 sky130_fd_sc_hd__xnor2_1 _5782_ (.A(_2298_),
    .B(_1624_),
    .Y(_2449_));
 sky130_fd_sc_hd__xnor2_1 _5783_ (.A(_2301_),
    .B(_1610_),
    .Y(_2452_));
 sky130_fd_sc_hd__nor2_1 _5784_ (.A(_2306_),
    .B(_1623_),
    .Y(_1625_));
 sky130_fd_sc_hd__xnor2_1 _5785_ (.A(_2304_),
    .B(_1625_),
    .Y(_2455_));
 sky130_fd_sc_hd__xnor2_1 _5786_ (.A(_2307_),
    .B(_1608_),
    .Y(_2458_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(_0142_),
    .B(_0143_),
    .Y(_1626_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(_2310_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__nor2_1 _5789_ (.A(_0144_),
    .B(_1627_),
    .Y(_2461_));
 sky130_fd_sc_hd__xor2_1 _5790_ (.A(_2108_),
    .B(_2313_),
    .X(_2464_));
 sky130_fd_sc_hd__nor3b_1 _5791_ (.A(_2412_),
    .B(_2416_),
    .C_N(_2329_),
    .Y(_1628_));
 sky130_fd_sc_hd__nor2_1 _5792_ (.A(net2),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__xor2_1 _5793_ (.A(_2408_),
    .B(_1629_),
    .X(_2477_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(net9),
    .B(_0764_),
    .Y(_1630_));
 sky130_fd_sc_hd__xnor2_1 _5795_ (.A(_2626_),
    .B(_1630_),
    .Y(_2485_));
 sky130_fd_sc_hd__xor2_1 _5796_ (.A(_2326_),
    .B(_2114_),
    .X(_2488_));
 sky130_fd_sc_hd__inv_1 _5797_ (.A(net33),
    .Y(_2509_));
 sky130_fd_sc_hd__inv_1 _5798_ (.A(net32),
    .Y(_2517_));
 sky130_fd_sc_hd__o31ai_1 _5799_ (.A1(_0682_),
    .A2(_0683_),
    .A3(_1596_),
    .B1(_0125_),
    .Y(_1631_));
 sky130_fd_sc_hd__xnor2_1 _5800_ (.A(_2574_),
    .B(_1631_),
    .Y(_2529_));
 sky130_fd_sc_hd__inv_1 _5801_ (.A(net35),
    .Y(_2541_));
 sky130_fd_sc_hd__inv_1 _5802_ (.A(net34),
    .Y(_2549_));
 sky130_fd_sc_hd__a31o_1 _5803_ (.A1(_2232_),
    .A2(_0684_),
    .A3(_1595_),
    .B1(net16),
    .X(_1632_));
 sky130_fd_sc_hd__xnor2_1 _5804_ (.A(_2562_),
    .B(_1632_),
    .Y(_2577_));
 sky130_fd_sc_hd__nor4_1 _5805_ (.A(_2760_),
    .B(_2728_),
    .C(_2732_),
    .D(_0794_),
    .Y(_1633_));
 sky130_fd_sc_hd__nor2_1 _5806_ (.A(net2),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__xor2_1 _5807_ (.A(_2764_),
    .B(_1634_),
    .X(_2585_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(_2728_),
    .B(_2732_),
    .Y(_1635_));
 sky130_fd_sc_hd__nor2_1 _5809_ (.A(_2404_),
    .B(_2408_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_1628_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__nor3_1 _5811_ (.A(_2534_),
    .B(_2538_),
    .C(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a21oi_1 _5812_ (.A1(_1635_),
    .A2(_1638_),
    .B1(_0159_),
    .Y(_1639_));
 sky130_fd_sc_hd__xor2_1 _5813_ (.A(_2760_),
    .B(_1639_),
    .X(_2589_));
 sky130_fd_sc_hd__o21ai_1 _5814_ (.A1(_2732_),
    .A2(_0794_),
    .B1(net18),
    .Y(_1640_));
 sky130_fd_sc_hd__xnor2_1 _5815_ (.A(_2728_),
    .B(_1640_),
    .Y(_2593_));
 sky130_fd_sc_hd__nor2_1 _5816_ (.A(net2),
    .B(_1638_),
    .Y(_1641_));
 sky130_fd_sc_hd__xor2_1 _5817_ (.A(_2732_),
    .B(_1641_),
    .X(_2597_));
 sky130_fd_sc_hd__o31ai_2 _5818_ (.A1(_2404_),
    .A2(_2538_),
    .A3(_0793_),
    .B1(_0295_),
    .Y(_1642_));
 sky130_fd_sc_hd__xnor2_1 _5819_ (.A(_2534_),
    .B(_1642_),
    .Y(_2601_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(net23),
    .B(_1637_),
    .Y(_1643_));
 sky130_fd_sc_hd__xnor2_1 _5821_ (.A(_2538_),
    .B(_1643_),
    .Y(_2605_));
 sky130_fd_sc_hd__nand2_1 _5822_ (.A(net23),
    .B(_0793_),
    .Y(_1644_));
 sky130_fd_sc_hd__xnor2_1 _5823_ (.A(_2404_),
    .B(_1644_),
    .Y(_2609_));
 sky130_fd_sc_hd__inv_1 _5824_ (.A(_2445_),
    .Y(_1645_));
 sky130_fd_sc_hd__inv_1 _5825_ (.A(_2125_),
    .Y(_1646_));
 sky130_fd_sc_hd__a21oi_1 _5826_ (.A1(_1646_),
    .A2(_2470_),
    .B1(_2469_),
    .Y(_1647_));
 sky130_fd_sc_hd__o21bai_1 _5827_ (.A1(_0331_),
    .A2(_1647_),
    .B1_N(_2467_),
    .Y(_1648_));
 sky130_fd_sc_hd__a21oi_1 _5828_ (.A1(_2466_),
    .A2(_1648_),
    .B1(_2465_),
    .Y(_1649_));
 sky130_fd_sc_hd__o21bai_1 _5829_ (.A1(_0330_),
    .A2(_1649_),
    .B1_N(_2462_),
    .Y(_1650_));
 sky130_fd_sc_hd__a21o_1 _5830_ (.A1(_2460_),
    .A2(_1650_),
    .B1(_2459_),
    .X(_1651_));
 sky130_fd_sc_hd__a21o_1 _5831_ (.A1(_2457_),
    .A2(_1651_),
    .B1(_2456_),
    .X(_1652_));
 sky130_fd_sc_hd__a21o_1 _5832_ (.A1(_2454_),
    .A2(_1652_),
    .B1(_2453_),
    .X(_1653_));
 sky130_fd_sc_hd__a21o_1 _5833_ (.A1(_2451_),
    .A2(_1653_),
    .B1(_2450_),
    .X(_1654_));
 sky130_fd_sc_hd__a21oi_1 _5834_ (.A1(_2448_),
    .A2(_1654_),
    .B1(_2447_),
    .Y(_1655_));
 sky130_fd_sc_hd__o21bai_1 _5835_ (.A1(_1645_),
    .A2(_1655_),
    .B1_N(_2444_),
    .Y(_1656_));
 sky130_fd_sc_hd__a21o_1 _5836_ (.A1(_2441_),
    .A2(_1656_),
    .B1(_2440_),
    .X(_1657_));
 sky130_fd_sc_hd__a21oi_1 _5837_ (.A1(_2438_),
    .A2(_1657_),
    .B1(_2437_),
    .Y(_1658_));
 sky130_fd_sc_hd__xnor2_1 _5838_ (.A(_2435_),
    .B(_1658_),
    .Y(_2651_));
 sky130_fd_sc_hd__o21bai_1 _5839_ (.A1(_1645_),
    .A2(_0342_),
    .B1_N(_2444_),
    .Y(_1659_));
 sky130_fd_sc_hd__a21oi_1 _5840_ (.A1(_2441_),
    .A2(_1659_),
    .B1(_2440_),
    .Y(_1660_));
 sky130_fd_sc_hd__xnor2_1 _5841_ (.A(_2438_),
    .B(_1660_),
    .Y(_2655_));
 sky130_fd_sc_hd__xor2_1 _5842_ (.A(_2441_),
    .B(_1656_),
    .X(_2658_));
 sky130_fd_sc_hd__xnor2_1 _5843_ (.A(_2445_),
    .B(_0342_),
    .Y(_2661_));
 sky130_fd_sc_hd__xor2_1 _5844_ (.A(_2448_),
    .B(_1654_),
    .X(_2664_));
 sky130_fd_sc_hd__nand2b_1 _5845_ (.A_N(_2453_),
    .B(_0338_),
    .Y(_1661_));
 sky130_fd_sc_hd__xor2_1 _5846_ (.A(_2451_),
    .B(_1661_),
    .X(_2668_));
 sky130_fd_sc_hd__xor2_1 _5847_ (.A(_2454_),
    .B(_1652_),
    .X(_2671_));
 sky130_fd_sc_hd__a21oi_1 _5848_ (.A1(_2460_),
    .A2(_0336_),
    .B1(_2459_),
    .Y(_1662_));
 sky130_fd_sc_hd__xnor2_1 _5849_ (.A(_2457_),
    .B(_1662_),
    .Y(_2674_));
 sky130_fd_sc_hd__xor2_1 _5850_ (.A(_2460_),
    .B(_1650_),
    .X(_2677_));
 sky130_fd_sc_hd__xnor2_1 _5851_ (.A(_2463_),
    .B(_0335_),
    .Y(_2680_));
 sky130_fd_sc_hd__xor2_1 _5852_ (.A(_2466_),
    .B(_1648_),
    .X(_2683_));
 sky130_fd_sc_hd__xnor2_1 _5853_ (.A(_2468_),
    .B(_0333_),
    .Y(_2686_));
 sky130_fd_sc_hd__xnor2_1 _5854_ (.A(_2125_),
    .B(_2470_),
    .Y(_2689_));
 sky130_fd_sc_hd__inv_1 _5855_ (.A(_2126_),
    .Y(_2692_));
 sky130_fd_sc_hd__o31ai_1 _5856_ (.A1(_2622_),
    .A2(_2626_),
    .A3(_0764_),
    .B1(_0578_),
    .Y(_1663_));
 sky130_fd_sc_hd__xnor2_1 _5857_ (.A(_2618_),
    .B(_1663_),
    .Y(_2695_));
 sky130_fd_sc_hd__nand2b_1 _5858_ (.A_N(_2822_),
    .B(_2716_),
    .Y(_1664_));
 sky130_fd_sc_hd__o21ai_0 _5859_ (.A1(_2818_),
    .A2(_1664_),
    .B1(_0816_),
    .Y(_1665_));
 sky130_fd_sc_hd__xnor2_1 _5860_ (.A(_2814_),
    .B(_1665_),
    .Y(_2703_));
 sky130_fd_sc_hd__xnor2_1 _5861_ (.A(_2487_),
    .B(_0636_),
    .Y(_2706_));
 sky130_fd_sc_hd__xor2_1 _5862_ (.A(_2129_),
    .B(_2491_),
    .X(_2710_));
 sky130_fd_sc_hd__or2b_1 _5863_ (.A(_2562_),
    .B_N(_0684_),
    .X(_1666_));
 sky130_fd_sc_hd__o21ai_1 _5864_ (.A1(_1666_),
    .A2(_0688_),
    .B1(net4),
    .Y(_1667_));
 sky130_fd_sc_hd__xnor2_1 _5865_ (.A(_2558_),
    .B(_1667_),
    .Y(_2723_));
 sky130_fd_sc_hd__o31ai_1 _5866_ (.A1(_2558_),
    .A2(_1666_),
    .A3(_1596_),
    .B1(_0125_),
    .Y(_1668_));
 sky130_fd_sc_hd__xnor2_1 _5867_ (.A(_0703_),
    .B(_1668_),
    .Y(_2735_));
 sky130_fd_sc_hd__xnor2_1 _5868_ (.A(_0782_),
    .B(_0796_),
    .Y(_2743_));
 sky130_fd_sc_hd__nor2_1 _5869_ (.A(_2944_),
    .B(_2928_),
    .Y(_1669_));
 sky130_fd_sc_hd__nor2_1 _5870_ (.A(_2630_),
    .B(_2626_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_2494_),
    .B(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__nor3_1 _5872_ (.A(_2622_),
    .B(_2618_),
    .C(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__nor2_1 _5873_ (.A(_2614_),
    .B(_2752_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _5874_ (.A(_1672_),
    .B(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__nor3_1 _5875_ (.A(_2748_),
    .B(_2932_),
    .C(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_1669_),
    .B(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _5877_ (.A(_0578_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__o31ai_1 _5878_ (.A1(_0783_),
    .A2(_0784_),
    .A3(_1677_),
    .B1(_0786_),
    .Y(_2767_));
 sky130_fd_sc_hd__nor2_1 _5879_ (.A(_0783_),
    .B(_0784_),
    .Y(_1678_));
 sky130_fd_sc_hd__xor2_1 _5880_ (.A(_1678_),
    .B(_1677_),
    .X(_2771_));
 sky130_fd_sc_hd__nor2_1 _5881_ (.A(_2665_),
    .B(_1675_),
    .Y(_1679_));
 sky130_fd_sc_hd__xor2_1 _5882_ (.A(_2928_),
    .B(_1679_),
    .X(_2777_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(net9),
    .B(_0767_),
    .Y(_1680_));
 sky130_fd_sc_hd__xnor2_1 _5884_ (.A(_2932_),
    .B(_1680_),
    .Y(_2781_));
 sky130_fd_sc_hd__nand2_1 _5885_ (.A(net9),
    .B(_1674_),
    .Y(_1681_));
 sky130_fd_sc_hd__xnor2_1 _5886_ (.A(_2748_),
    .B(_1681_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand2_1 _5887_ (.A(net9),
    .B(_0766_),
    .Y(_1682_));
 sky130_fd_sc_hd__xnor2_1 _5888_ (.A(_2752_),
    .B(_1682_),
    .Y(_2789_));
 sky130_fd_sc_hd__nor2_1 _5889_ (.A(_2665_),
    .B(_1672_),
    .Y(_1683_));
 sky130_fd_sc_hd__xnor2_1 _5890_ (.A(_0438_),
    .B(_1683_),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(_0785_),
    .B(_0786_),
    .Y(_2797_));
 sky130_fd_sc_hd__o31ai_1 _5892_ (.A1(_2928_),
    .A2(_2932_),
    .A3(_0767_),
    .B1(_0578_),
    .Y(_1684_));
 sky130_fd_sc_hd__xnor2_1 _5893_ (.A(_2944_),
    .B(_1684_),
    .Y(_2801_));
 sky130_fd_sc_hd__inv_1 _5894_ (.A(_2337_),
    .Y(_2131_));
 sky130_fd_sc_hd__nor2_1 _5895_ (.A(_2476_),
    .B(_0348_),
    .Y(_1685_));
 sky130_fd_sc_hd__a21oi_1 _5896_ (.A1(_0138_),
    .A2(_2476_),
    .B1(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a21oi_1 _5897_ (.A1(_2691_),
    .A2(_1686_),
    .B1(_2690_),
    .Y(_1687_));
 sky130_fd_sc_hd__nor2b_1 _5898_ (.A(_1687_),
    .B_N(_2688_),
    .Y(_1688_));
 sky130_fd_sc_hd__o21ai_0 _5899_ (.A1(_2687_),
    .A2(_1688_),
    .B1(_2685_),
    .Y(_1689_));
 sky130_fd_sc_hd__a21boi_0 _5900_ (.A1(_0612_),
    .A2(_1689_),
    .B1_N(_2682_),
    .Y(_1690_));
 sky130_fd_sc_hd__o21a_1 _5901_ (.A1(_2681_),
    .A2(_1690_),
    .B1(_2679_),
    .X(_1691_));
 sky130_fd_sc_hd__o21a_1 _5902_ (.A1(_2678_),
    .A2(_1691_),
    .B1(_2676_),
    .X(_1692_));
 sky130_fd_sc_hd__o21a_1 _5903_ (.A1(_2675_),
    .A2(_1692_),
    .B1(_2673_),
    .X(_1693_));
 sky130_fd_sc_hd__o21a_1 _5904_ (.A1(_2672_),
    .A2(_1693_),
    .B1(_2670_),
    .X(_1694_));
 sky130_fd_sc_hd__o21a_1 _5905_ (.A1(_2669_),
    .A2(_1694_),
    .B1(_2667_),
    .X(_1695_));
 sky130_fd_sc_hd__o21a_1 _5906_ (.A1(_2666_),
    .A2(_1695_),
    .B1(_2663_),
    .X(_1696_));
 sky130_fd_sc_hd__o21ai_0 _5907_ (.A1(_2662_),
    .A2(_1696_),
    .B1(_2660_),
    .Y(_1697_));
 sky130_fd_sc_hd__nand2b_1 _5908_ (.A_N(_2659_),
    .B(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__a21oi_1 _5909_ (.A1(_2657_),
    .A2(_1698_),
    .B1(_2656_),
    .Y(_1699_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(_2654_),
    .B(_1699_),
    .Y(_2851_));
 sky130_fd_sc_hd__a21oi_1 _5911_ (.A1(_2660_),
    .A2(_0626_),
    .B1(_2659_),
    .Y(_1700_));
 sky130_fd_sc_hd__xnor2_1 _5912_ (.A(_2657_),
    .B(_1700_),
    .Y(_2855_));
 sky130_fd_sc_hd__nor2_1 _5913_ (.A(_2662_),
    .B(_1696_),
    .Y(_1701_));
 sky130_fd_sc_hd__xnor2_1 _5914_ (.A(_2660_),
    .B(_1701_),
    .Y(_2858_));
 sky130_fd_sc_hd__xor2_1 _5915_ (.A(_2663_),
    .B(_0625_),
    .X(_2861_));
 sky130_fd_sc_hd__nor3_1 _5916_ (.A(_2667_),
    .B(_2669_),
    .C(_1694_),
    .Y(_1702_));
 sky130_fd_sc_hd__nor2_1 _5917_ (.A(_1695_),
    .B(_1702_),
    .Y(_2864_));
 sky130_fd_sc_hd__nor2_1 _5918_ (.A(_0621_),
    .B(_0622_),
    .Y(_1703_));
 sky130_fd_sc_hd__xnor2_1 _5919_ (.A(_2670_),
    .B(_1703_),
    .Y(_2867_));
 sky130_fd_sc_hd__nor3_1 _5920_ (.A(_2673_),
    .B(_2675_),
    .C(_1692_),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _5921_ (.A(_1693_),
    .B(_1704_),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _5922_ (.A(_0611_),
    .B(_0619_),
    .Y(_1705_));
 sky130_fd_sc_hd__xor2_1 _5923_ (.A(_2676_),
    .B(_1705_),
    .X(_2874_));
 sky130_fd_sc_hd__nor3_1 _5924_ (.A(_2679_),
    .B(_2681_),
    .C(_1690_),
    .Y(_1706_));
 sky130_fd_sc_hd__nor2_1 _5925_ (.A(_1691_),
    .B(_1706_),
    .Y(_2877_));
 sky130_fd_sc_hd__nand2_1 _5926_ (.A(_0612_),
    .B(_0617_),
    .Y(_1707_));
 sky130_fd_sc_hd__nor2_1 _5927_ (.A(_2682_),
    .B(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__nor2_1 _5928_ (.A(_0618_),
    .B(_1708_),
    .Y(_2880_));
 sky130_fd_sc_hd__nor2_1 _5929_ (.A(_2687_),
    .B(_1688_),
    .Y(_1709_));
 sky130_fd_sc_hd__xnor2_1 _5930_ (.A(_2685_),
    .B(_1709_),
    .Y(_2883_));
 sky130_fd_sc_hd__nand2_1 _5931_ (.A(_0613_),
    .B(_0615_),
    .Y(_1710_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(_2688_),
    .B(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__nor2_1 _5933_ (.A(_0616_),
    .B(_1711_),
    .Y(_2886_));
 sky130_fd_sc_hd__xor2_1 _5934_ (.A(_2691_),
    .B(_1686_),
    .X(_2889_));
 sky130_fd_sc_hd__xnor2_1 _5935_ (.A(_0138_),
    .B(_2694_),
    .Y(_2892_));
 sky130_fd_sc_hd__or4_1 _5936_ (.A(_2848_),
    .B(_2818_),
    .C(_2814_),
    .D(_1664_),
    .X(_1712_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(net12),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__xnor2_1 _5938_ (.A(_2810_),
    .B(_1713_),
    .Y(_2895_));
 sky130_fd_sc_hd__o21ai_0 _5939_ (.A1(_1101_),
    .A2(_1102_),
    .B1(_0972_),
    .Y(_1714_));
 sky130_fd_sc_hd__xnor2_1 _5940_ (.A(_2986_),
    .B(_1714_),
    .Y(_2903_));
 sky130_fd_sc_hd__xnor2_1 _5941_ (.A(_2705_),
    .B(_0877_),
    .Y(_2906_));
 sky130_fd_sc_hd__xnor2_1 _5942_ (.A(_2709_),
    .B(_0644_),
    .Y(_2910_));
 sky130_fd_sc_hd__xor2_1 _5943_ (.A(_2713_),
    .B(_2138_),
    .X(_2914_));
 sky130_fd_sc_hd__inv_1 _5944_ (.A(_2940_),
    .Y(_1715_));
 sky130_fd_sc_hd__nor3_1 _5945_ (.A(_2806_),
    .B(_2810_),
    .C(_1712_),
    .Y(_1716_));
 sky130_fd_sc_hd__nand3_1 _5946_ (.A(_0908_),
    .B(_1715_),
    .C(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__or2_0 _5947_ (.A(_0950_),
    .B(_0951_),
    .X(_1718_));
 sky130_fd_sc_hd__o211ai_1 _5948_ (.A1(_3117_),
    .A2(_1717_),
    .B1(_1718_),
    .C1(net12),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(_0952_),
    .B(_1719_),
    .Y(_2947_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_0952_),
    .B(_1719_),
    .Y(_2951_));
 sky130_fd_sc_hd__nand2_1 _5951_ (.A(net12),
    .B(_1717_),
    .Y(_1720_));
 sky130_fd_sc_hd__xnor2_1 _5952_ (.A(_3117_),
    .B(_1720_),
    .Y(_2957_));
 sky130_fd_sc_hd__nor2_1 _5953_ (.A(net1),
    .B(_0956_),
    .Y(_1721_));
 sky130_fd_sc_hd__xnor2_1 _5954_ (.A(_0908_),
    .B(_1721_),
    .Y(_2961_));
 sky130_fd_sc_hd__nor2_1 _5955_ (.A(net1),
    .B(_1716_),
    .Y(_1722_));
 sky130_fd_sc_hd__xnor2_1 _5956_ (.A(_1715_),
    .B(_1722_),
    .Y(_2965_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(net12),
    .B(_0955_),
    .Y(_1723_));
 sky130_fd_sc_hd__xnor2_1 _5958_ (.A(_2806_),
    .B(_1723_),
    .Y(_2969_));
 sky130_fd_sc_hd__xnor2_1 _5959_ (.A(_1718_),
    .B(_0957_),
    .Y(_2977_));
 sky130_fd_sc_hd__inv_1 _5960_ (.A(_2144_),
    .Y(_2154_));
 sky130_fd_sc_hd__inv_1 _5961_ (.A(_2872_),
    .Y(_1724_));
 sky130_fd_sc_hd__inv_1 _5962_ (.A(_2878_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_0138_),
    .B(_2694_),
    .Y(_1726_));
 sky130_fd_sc_hd__o21ai_1 _5964_ (.A1(_2694_),
    .A2(net13),
    .B1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__a21oi_1 _5965_ (.A1(_2891_),
    .A2(_1727_),
    .B1(_2890_),
    .Y(_1728_));
 sky130_fd_sc_hd__o21ai_1 _5966_ (.A1(_0857_),
    .A2(_1728_),
    .B1(_0860_),
    .Y(_1729_));
 sky130_fd_sc_hd__a21oi_1 _5967_ (.A1(_2885_),
    .A2(_1729_),
    .B1(_2884_),
    .Y(_1730_));
 sky130_fd_sc_hd__nor2_1 _5968_ (.A(_0856_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__o21ai_0 _5969_ (.A1(_2881_),
    .A2(_1731_),
    .B1(_2879_),
    .Y(_1732_));
 sky130_fd_sc_hd__a21oi_1 _5970_ (.A1(_1725_),
    .A2(_1732_),
    .B1(_0855_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21ai_0 _5971_ (.A1(_2875_),
    .A2(_1733_),
    .B1(_2873_),
    .Y(_1734_));
 sky130_fd_sc_hd__a21oi_1 _5972_ (.A1(_1724_),
    .A2(_1734_),
    .B1(_0854_),
    .Y(_1735_));
 sky130_fd_sc_hd__o21a_1 _5973_ (.A1(_2869_),
    .A2(_1735_),
    .B1(_2866_),
    .X(_1736_));
 sky130_fd_sc_hd__o21ai_0 _5974_ (.A1(_2865_),
    .A2(_1736_),
    .B1(_2863_),
    .Y(_1737_));
 sky130_fd_sc_hd__nand2b_1 _5975_ (.A_N(_2862_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__a21o_1 _5976_ (.A1(_2860_),
    .A2(_1738_),
    .B1(_2859_),
    .X(_1739_));
 sky130_fd_sc_hd__a21oi_1 _5977_ (.A1(_2857_),
    .A2(_1739_),
    .B1(_2856_),
    .Y(_1740_));
 sky130_fd_sc_hd__xnor2_1 _5978_ (.A(_2854_),
    .B(_1740_),
    .Y(_3037_));
 sky130_fd_sc_hd__xnor2_1 _5979_ (.A(_2857_),
    .B(_0870_),
    .Y(_3041_));
 sky130_fd_sc_hd__xor2_1 _5980_ (.A(_2860_),
    .B(_1738_),
    .X(_3044_));
 sky130_fd_sc_hd__xnor2_1 _5981_ (.A(_2863_),
    .B(_0868_),
    .Y(_3047_));
 sky130_fd_sc_hd__nor2_1 _5982_ (.A(_2869_),
    .B(_1735_),
    .Y(_1741_));
 sky130_fd_sc_hd__xnor2_1 _5983_ (.A(_2866_),
    .B(_1741_),
    .Y(_3050_));
 sky130_fd_sc_hd__xnor2_1 _5984_ (.A(_2870_),
    .B(_0866_),
    .Y(_3053_));
 sky130_fd_sc_hd__nor2_1 _5985_ (.A(_2875_),
    .B(_1733_),
    .Y(_1742_));
 sky130_fd_sc_hd__xnor2_1 _5986_ (.A(_2873_),
    .B(_1742_),
    .Y(_3056_));
 sky130_fd_sc_hd__xnor2_1 _5987_ (.A(_2876_),
    .B(_0864_),
    .Y(_3060_));
 sky130_fd_sc_hd__nor2_1 _5988_ (.A(_2881_),
    .B(_1731_),
    .Y(_1743_));
 sky130_fd_sc_hd__xnor2_1 _5989_ (.A(_2879_),
    .B(_1743_),
    .Y(_3063_));
 sky130_fd_sc_hd__xnor2_1 _5990_ (.A(_2882_),
    .B(_0862_),
    .Y(_3066_));
 sky130_fd_sc_hd__xor2_1 _5991_ (.A(_2885_),
    .B(_1729_),
    .X(_3069_));
 sky130_fd_sc_hd__xnor2_1 _5992_ (.A(_2888_),
    .B(_0859_),
    .Y(_3072_));
 sky130_fd_sc_hd__xor2_1 _5993_ (.A(_2891_),
    .B(_1727_),
    .X(_3075_));
 sky130_fd_sc_hd__xor2_2 _5994_ (.A(_0138_),
    .B(_2894_),
    .X(_3078_));
 sky130_fd_sc_hd__nand2_1 _5995_ (.A(net24),
    .B(_1103_),
    .Y(_1744_));
 sky130_fd_sc_hd__xnor2_1 _5996_ (.A(_3029_),
    .B(_1744_),
    .Y(_3081_));
 sky130_fd_sc_hd__a21oi_1 _5997_ (.A1(_1235_),
    .A2(_1237_),
    .B1(net25),
    .Y(_1745_));
 sky130_fd_sc_hd__xor2_1 _5998_ (.A(_3197_),
    .B(_1745_),
    .X(_3085_));
 sky130_fd_sc_hd__nor2b_2 _5999_ (.A(_3163_),
    .B_N(_3110_),
    .Y(_1746_));
 sky130_fd_sc_hd__a21oi_1 _6000_ (.A1(_1236_),
    .A2(_1746_),
    .B1(_1049_),
    .Y(_1747_));
 sky130_fd_sc_hd__xor2_1 _6001_ (.A(_3201_),
    .B(_1747_),
    .X(_3089_));
 sky130_fd_sc_hd__xnor2_2 _6002_ (.A(_2905_),
    .B(_1054_),
    .Y(_3092_));
 sky130_fd_sc_hd__xnor2_2 _6003_ (.A(_2909_),
    .B(_0894_),
    .Y(_3096_));
 sky130_fd_sc_hd__xnor2_2 _6004_ (.A(_2913_),
    .B(_1052_),
    .Y(_3100_));
 sky130_fd_sc_hd__xor2_2 _6005_ (.A(_2148_),
    .B(_2917_),
    .X(_3104_));
 sky130_fd_sc_hd__or2_1 _6006_ (.A(_1098_),
    .B(_1099_),
    .X(_1748_));
 sky130_fd_sc_hd__nand2b_1 _6007_ (.A_N(_3000_),
    .B(_2920_),
    .Y(_1749_));
 sky130_fd_sc_hd__nor3_1 _6008_ (.A(_2986_),
    .B(_1102_),
    .C(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__nor2_1 _6009_ (.A(_3034_),
    .B(_3029_),
    .Y(_1751_));
 sky130_fd_sc_hd__nand2_1 _6010_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__o31ai_2 _6011_ (.A1(_2981_),
    .A2(_3121_),
    .A3(_1752_),
    .B1(net17),
    .Y(_1753_));
 sky130_fd_sc_hd__o21bai_1 _6012_ (.A1(_1748_),
    .A2(_1753_),
    .B1_N(_1106_),
    .Y(_3125_));
 sky130_fd_sc_hd__xnor2_1 _6013_ (.A(_1748_),
    .B(_1753_),
    .Y(_3137_));
 sky130_fd_sc_hd__o31ai_1 _6014_ (.A1(_2981_),
    .A2(_3029_),
    .A3(_1103_),
    .B1(net24),
    .Y(_1754_));
 sky130_fd_sc_hd__xnor2_1 _6015_ (.A(_3121_),
    .B(_1754_),
    .Y(_3141_));
 sky130_fd_sc_hd__nand2_1 _6016_ (.A(net24),
    .B(_1752_),
    .Y(_1755_));
 sky130_fd_sc_hd__xnor2_1 _6017_ (.A(_2981_),
    .B(_1755_),
    .Y(_3145_));
 sky130_fd_sc_hd__o21bai_1 _6018_ (.A1(_1748_),
    .A2(_1753_),
    .B1_N(_1106_),
    .Y(_3133_));
 sky130_fd_sc_hd__or2_0 _6019_ (.A(_1105_),
    .B(_1106_),
    .X(_3151_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_0991_),
    .B(_0993_),
    .Y(_1756_));
 sky130_fd_sc_hd__nor2_1 _6021_ (.A(_3018_),
    .B(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__nor2_1 _6022_ (.A(_0994_),
    .B(_1757_),
    .Y(_3183_));
 sky130_fd_sc_hd__inv_1 _6023_ (.A(_2153_),
    .Y(_2160_));
 sky130_fd_sc_hd__mux2i_2 _6024_ (.A0(_3057_),
    .A1(net28),
    .S(_2894_),
    .Y(_1758_));
 sky130_fd_sc_hd__a21oi_1 _6025_ (.A1(_3077_),
    .A2(_1758_),
    .B1(_3076_),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2b_1 _6026_ (.A(_1759_),
    .B_N(_3074_),
    .Y(_1760_));
 sky130_fd_sc_hd__o21ai_0 _6027_ (.A1(_3073_),
    .A2(_1760_),
    .B1(_3071_),
    .Y(_1761_));
 sky130_fd_sc_hd__a21boi_0 _6028_ (.A1(_1032_),
    .A2(_1761_),
    .B1_N(_3068_),
    .Y(_1762_));
 sky130_fd_sc_hd__nor2_1 _6029_ (.A(_3067_),
    .B(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hd__xnor2_1 _6030_ (.A(_3065_),
    .B(_1763_),
    .Y(_3239_));
 sky130_fd_sc_hd__xnor2_1 _6031_ (.A(net28),
    .B(_3080_),
    .Y(_3254_));
 sky130_fd_sc_hd__xnor2_1 _6032_ (.A(_3091_),
    .B(_1193_),
    .Y(_3265_));
 sky130_fd_sc_hd__o21ai_0 _6033_ (.A1(_3368_),
    .A2(_1459_),
    .B1(net20),
    .Y(_1764_));
 sky130_fd_sc_hd__xnor2_1 _6034_ (.A(_3365_),
    .B(_1764_),
    .Y(_3269_));
 sky130_fd_sc_hd__nor3b_1 _6035_ (.A(_3324_),
    .B(_3372_),
    .C_N(_3287_),
    .Y(_1765_));
 sky130_fd_sc_hd__nor2_1 _6036_ (.A(_3405_),
    .B(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__xor2_1 _6037_ (.A(_3368_),
    .B(_1766_),
    .X(_3273_));
 sky130_fd_sc_hd__nor2_1 _6038_ (.A(_1186_),
    .B(_1458_),
    .Y(_1767_));
 sky130_fd_sc_hd__xor2_1 _6039_ (.A(_3324_),
    .B(_1767_),
    .X(_3277_));
 sky130_fd_sc_hd__nor2_4 _6040_ (.A(_3405_),
    .B(_3287_),
    .Y(_1768_));
 sky130_fd_sc_hd__xor2_1 _6041_ (.A(_3372_),
    .B(_1768_),
    .X(_3281_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_3288_),
    .B(_3380_),
    .Y(_1769_));
 sky130_fd_sc_hd__o21ai_2 _6043_ (.A1(_3285_),
    .A2(_3380_),
    .B1(_1769_),
    .Y(_2167_));
 sky130_fd_sc_hd__xnor2_1 _6044_ (.A(_3174_),
    .B(_1145_),
    .Y(_3332_));
 sky130_fd_sc_hd__xor2_1 _6045_ (.A(_3178_),
    .B(_1157_),
    .X(_3338_));
 sky130_fd_sc_hd__xor2_1 _6046_ (.A(_3186_),
    .B(_1155_),
    .X(_3346_));
 sky130_fd_sc_hd__xor2_1 _6047_ (.A(_2163_),
    .B(_3190_),
    .X(_3350_));
 sky130_fd_sc_hd__nand2_4 _6048_ (.A(_1462_),
    .B(_1463_),
    .Y(_1770_));
 sky130_fd_sc_hd__nor2b_1 _6049_ (.A(_1460_),
    .B_N(_1765_),
    .Y(_1771_));
 sky130_fd_sc_hd__nor2_1 _6050_ (.A(_3321_),
    .B(_3361_),
    .Y(_1772_));
 sky130_fd_sc_hd__a21oi_2 _6051_ (.A1(_1771_),
    .A2(_1772_),
    .B1(_1186_),
    .Y(_1773_));
 sky130_fd_sc_hd__xor2_2 _6052_ (.A(_1773_),
    .B(_1770_),
    .X(_3261_));
 sky130_fd_sc_hd__nand2_1 _6053_ (.A(net7),
    .B(_1461_),
    .Y(_1774_));
 sky130_fd_sc_hd__xnor2_1 _6054_ (.A(_3321_),
    .B(_1774_),
    .Y(_3430_));
 sky130_fd_sc_hd__nor2_1 _6055_ (.A(_1319_),
    .B(_1358_),
    .Y(_1775_));
 sky130_fd_sc_hd__xor2_1 _6056_ (.A(_3649_),
    .B(_1775_),
    .X(_3444_));
 sky130_fd_sc_hd__xnor2_1 _6057_ (.A(_3280_),
    .B(_1333_),
    .Y(_3448_));
 sky130_fd_sc_hd__o21ai_0 _6058_ (.A1(_3620_),
    .A2(_1356_),
    .B1(_3489_),
    .Y(_1776_));
 sky130_fd_sc_hd__xnor2_1 _6059_ (.A(_3633_),
    .B(_1776_),
    .Y(_3452_));
 sky130_fd_sc_hd__xnor2_2 _6060_ (.A(_3432_),
    .B(_1337_),
    .Y(_3473_));
 sky130_fd_sc_hd__nor2_1 _6061_ (.A(_1319_),
    .B(_1360_),
    .Y(_1777_));
 sky130_fd_sc_hd__xor2_1 _6062_ (.A(_3665_),
    .B(_1777_),
    .X(_3477_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_1319_),
    .B(_1359_),
    .Y(_1778_));
 sky130_fd_sc_hd__xor2_1 _6064_ (.A(_3657_),
    .B(_1778_),
    .X(_3481_));
 sky130_fd_sc_hd__inv_1 _6065_ (.A(net214),
    .Y(_3485_));
 sky130_fd_sc_hd__inv_1 _6066_ (.A(_3401_),
    .Y(_1779_));
 sky130_fd_sc_hd__inv_1 _6067_ (.A(_3408_),
    .Y(_1780_));
 sky130_fd_sc_hd__a211oi_1 _6068_ (.A1(_3216_),
    .A2(_1184_),
    .B1(_3256_),
    .C1(_3215_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _6069_ (.A(net28),
    .B(_3256_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_3420_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__o21bai_1 _6071_ (.A1(_1781_),
    .A2(_1783_),
    .B1_N(_3419_),
    .Y(_1784_));
 sky130_fd_sc_hd__a21o_1 _6072_ (.A1(_3417_),
    .A2(_1784_),
    .B1(_3416_),
    .X(_1785_));
 sky130_fd_sc_hd__a21o_1 _6073_ (.A1(_3414_),
    .A2(_1785_),
    .B1(_3413_),
    .X(_1786_));
 sky130_fd_sc_hd__a21oi_1 _6074_ (.A1(_3411_),
    .A2(_1786_),
    .B1(_3410_),
    .Y(_1787_));
 sky130_fd_sc_hd__o21ai_0 _6075_ (.A1(_1780_),
    .A2(_1787_),
    .B1(_1297_),
    .Y(_1788_));
 sky130_fd_sc_hd__a21oi_1 _6076_ (.A1(_3404_),
    .A2(_1788_),
    .B1(_3403_),
    .Y(_1789_));
 sky130_fd_sc_hd__o21ai_0 _6077_ (.A1(_1779_),
    .A2(_1789_),
    .B1(_1296_),
    .Y(_1790_));
 sky130_fd_sc_hd__a21oi_1 _6078_ (.A1(_3398_),
    .A2(_1790_),
    .B1(_3397_),
    .Y(_1791_));
 sky130_fd_sc_hd__nor2b_1 _6079_ (.A(_1791_),
    .B_N(_3395_),
    .Y(_1792_));
 sky130_fd_sc_hd__o21ai_0 _6080_ (.A1(_3394_),
    .A2(_1792_),
    .B1(_3392_),
    .Y(_1793_));
 sky130_fd_sc_hd__nand2b_1 _6081_ (.A_N(_3391_),
    .B(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__xor2_1 _6082_ (.A(_3389_),
    .B(_1794_),
    .X(_3496_));
 sky130_fd_sc_hd__xor2_1 _6083_ (.A(_3392_),
    .B(_1310_),
    .X(_3499_));
 sky130_fd_sc_hd__xor2_1 _6084_ (.A(_3414_),
    .B(_1785_),
    .X(_3521_));
 sky130_fd_sc_hd__inv_1 _6085_ (.A(_2179_),
    .Y(_2185_));
 sky130_fd_sc_hd__nor2_2 _6086_ (.A(_3461_),
    .B(_3517_),
    .Y(_1795_));
 sky130_fd_sc_hd__xnor2_1 _6087_ (.A(_1795_),
    .B(_3469_),
    .Y(_3529_));
 sky130_fd_sc_hd__nor2_2 _6088_ (.A(_1397_),
    .B(_3487_),
    .Y(_1796_));
 sky130_fd_sc_hd__xnor2_1 _6089_ (.A(net137),
    .B(_1796_),
    .Y(_3541_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_3489_),
    .B(_1489_),
    .Y(_1797_));
 sky130_fd_sc_hd__xor2_1 _6091_ (.A(_3537_),
    .B(_1797_),
    .X(_3545_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_1431_),
    .B(_1433_),
    .Y(_3553_));
 sky130_fd_sc_hd__xor2_1 _6093_ (.A(_3548_),
    .B(net155),
    .X(_3557_));
 sky130_fd_sc_hd__nor2_1 _6094_ (.A(_3517_),
    .B(_1473_),
    .Y(_1798_));
 sky130_fd_sc_hd__xnor2_1 _6095_ (.A(_3554_),
    .B(_1798_),
    .Y(_3561_));
 sky130_fd_sc_hd__xor2_2 _6096_ (.A(_3564_),
    .B(net131),
    .X(_3573_));
 sky130_fd_sc_hd__xor2_2 _6097_ (.A(_3341_),
    .B(_1284_),
    .X(_3577_));
 sky130_fd_sc_hd__xor2_2 _6098_ (.A(_3580_),
    .B(_1497_),
    .X(_3589_));
 sky130_fd_sc_hd__xor2_2 _6099_ (.A(_3335_),
    .B(_1271_),
    .X(_3593_));
 sky130_fd_sc_hd__xor2_2 _6100_ (.A(_3596_),
    .B(net150),
    .X(_3601_));
 sky130_fd_sc_hd__nand2_4 _6101_ (.A(_3608_),
    .B(_3489_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand2_4 _6102_ (.A(_1556_),
    .B(_1799_),
    .Y(_3609_));
 sky130_fd_sc_hd__a31o_1 _6103_ (.A1(_1485_),
    .A2(_1486_),
    .A3(_1488_),
    .B1(_1504_),
    .X(_3613_));
 sky130_fd_sc_hd__nor2_1 _6104_ (.A(_3615_),
    .B(_1397_),
    .Y(_1800_));
 sky130_fd_sc_hd__nor2_1 _6105_ (.A(_1800_),
    .B(_1507_),
    .Y(_3616_));
 sky130_fd_sc_hd__xor2_2 _6106_ (.A(net213),
    .B(net151),
    .X(_3624_));
 sky130_fd_sc_hd__nand2_4 _6107_ (.A(_3675_),
    .B(_1555_),
    .Y(_1801_));
 sky130_fd_sc_hd__o21ai_4 _6108_ (.A1(_1555_),
    .A2(net238),
    .B1(_1801_),
    .Y(_2192_));
 sky130_fd_sc_hd__xor2_2 _6109_ (.A(_2189_),
    .B(_3455_),
    .X(_3689_));
 sky130_fd_sc_hd__xnor2_2 _6110_ (.A(_3451_),
    .B(_1345_),
    .Y(_3693_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_3674_),
    .B(_1535_),
    .Y(_1802_));
 sky130_fd_sc_hd__o21ai_0 _6112_ (.A1(_3653_),
    .A2(_1802_),
    .B1(_1555_),
    .Y(_1803_));
 sky130_fd_sc_hd__xnor2_1 _6113_ (.A(_3661_),
    .B(_1803_),
    .Y(_3697_));
 sky130_fd_sc_hd__nand4bb_4 _6114_ (.A_N(net153),
    .B_N(_1525_),
    .C(_1526_),
    .D(net191),
    .Y(_1804_));
 sky130_fd_sc_hd__o31ai_2 _6115_ (.A1(_3653_),
    .A2(_3661_),
    .A3(_1804_),
    .B1(_1555_),
    .Y(_1805_));
 sky130_fd_sc_hd__xnor2_1 _6116_ (.A(_3669_),
    .B(_1805_),
    .Y(_3701_));
 sky130_fd_sc_hd__xnor2_2 _6117_ (.A(_3480_),
    .B(_1367_),
    .Y(_3709_));
 sky130_fd_sc_hd__a21oi_2 _6118_ (.A1(net197),
    .A2(_1568_),
    .B1(_1398_),
    .Y(_1806_));
 sky130_fd_sc_hd__o21bai_1 _6119_ (.A1(_3715_),
    .A2(_1397_),
    .B1_N(_1806_),
    .Y(_3716_));
 sky130_fd_sc_hd__xnor2_2 _6120_ (.A(_3439_),
    .B(net161),
    .Y(_3720_));
 sky130_fd_sc_hd__nor4_2 _6121_ (.A(_3653_),
    .B(_3661_),
    .C(_3669_),
    .D(_1804_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand3_1 _6122_ (.A(_1555_),
    .B(net197),
    .C(_1568_),
    .Y(_1808_));
 sky130_fd_sc_hd__o21bai_1 _6123_ (.A1(_1807_),
    .A2(_1808_),
    .B1_N(_1806_),
    .Y(_3739_));
 sky130_fd_sc_hd__inv_1 _6124_ (.A(net46),
    .Y(_2197_));
 sky130_fd_sc_hd__inv_1 _6125_ (.A(net53),
    .Y(_2082_));
 sky130_fd_sc_hd__inv_1 _6126_ (.A(net55),
    .Y(_2212_));
 sky130_fd_sc_hd__inv_1 _6127_ (.A(net54),
    .Y(_2220_));
 sky130_fd_sc_hd__nor2_1 _6128_ (.A(_2232_),
    .B(net16),
    .Y(_1809_));
 sky130_fd_sc_hd__xnor2_1 _6129_ (.A(_0031_),
    .B(_1809_),
    .Y(_2228_));
 sky130_fd_sc_hd__inv_1 _6130_ (.A(net57),
    .Y(_2242_));
 sky130_fd_sc_hd__inv_1 _6131_ (.A(net56),
    .Y(_2250_));
 sky130_fd_sc_hd__inv_1 _6132_ (.A(net58),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _6133_ (.A(net23),
    .B(_0792_),
    .Y(_1810_));
 sky130_fd_sc_hd__xnor2_1 _6134_ (.A(_2412_),
    .B(_1810_),
    .Y(_2321_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_2330_),
    .B(net23),
    .Y(_1811_));
 sky130_fd_sc_hd__o21ai_1 _6136_ (.A1(_2328_),
    .A2(_2124_),
    .B1(_1811_),
    .Y(_2113_));
 sky130_fd_sc_hd__inv_1 _6137_ (.A(_2196_),
    .Y(_2334_));
 sky130_fd_sc_hd__inv_1 _6138_ (.A(net59),
    .Y(_2342_));
 sky130_fd_sc_hd__inv_1 _6139_ (.A(net60),
    .Y(_2350_));
 sky130_fd_sc_hd__inv_1 _6140_ (.A(net47),
    .Y(_2366_));
 sky130_fd_sc_hd__inv_1 _6141_ (.A(net61),
    .Y(_2374_));
 sky130_fd_sc_hd__o31ai_1 _6142_ (.A1(_2502_),
    .A2(_0682_),
    .A3(_0688_),
    .B1(_0125_),
    .Y(_1812_));
 sky130_fd_sc_hd__xnor2_1 _6143_ (.A(_2570_),
    .B(_1812_),
    .Y(_2380_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(net9),
    .B(_1671_),
    .Y(_1813_));
 sky130_fd_sc_hd__xnor2_1 _6145_ (.A(_2622_),
    .B(_1813_),
    .Y(_2482_));
 sky130_fd_sc_hd__nor2_1 _6146_ (.A(_2494_),
    .B(_2665_),
    .Y(_1814_));
 sky130_fd_sc_hd__xor2_1 _6147_ (.A(_2630_),
    .B(_1814_),
    .X(_2489_));
 sky130_fd_sc_hd__nand2_1 _6148_ (.A(_2495_),
    .B(net9),
    .Y(_1815_));
 sky130_fd_sc_hd__o21ai_1 _6149_ (.A1(_2493_),
    .A2(net9),
    .B1(_1815_),
    .Y(_2128_));
 sky130_fd_sc_hd__inv_1 _6150_ (.A(net49),
    .Y(_2512_));
 sky130_fd_sc_hd__inv_1 _6151_ (.A(net48),
    .Y(_2520_));
 sky130_fd_sc_hd__o41ai_1 _6152_ (.A1(_2574_),
    .A2(_0682_),
    .A3(_0683_),
    .A4(_0688_),
    .B1(_0115_),
    .Y(_1816_));
 sky130_fd_sc_hd__xnor2_1 _6153_ (.A(_2566_),
    .B(_1816_),
    .Y(_2526_));
 sky130_fd_sc_hd__inv_1 _6154_ (.A(net51),
    .Y(_2544_));
 sky130_fd_sc_hd__inv_1 _6155_ (.A(net50),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_0791_),
    .B(_1638_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _6157_ (.A(net23),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__xnor2_1 _6158_ (.A(_2756_),
    .B(_1818_),
    .Y(_2582_));
 sky130_fd_sc_hd__xnor2_1 _6159_ (.A(_2119_),
    .B(_2426_),
    .Y(_2642_));
 sky130_fd_sc_hd__inv_1 _6160_ (.A(_2120_),
    .Y(_2133_));
 sky130_fd_sc_hd__nand2_1 _6161_ (.A(net12),
    .B(_0954_),
    .Y(_1819_));
 sky130_fd_sc_hd__xnor2_1 _6162_ (.A(_2848_),
    .B(_1819_),
    .Y(_2700_));
 sky130_fd_sc_hd__nand2_1 _6163_ (.A(net12),
    .B(_0953_),
    .Y(_1820_));
 sky130_fd_sc_hd__xnor2_1 _6164_ (.A(_2818_),
    .B(_1820_),
    .Y(_2707_));
 sky130_fd_sc_hd__nor2_1 _6165_ (.A(_2716_),
    .B(net1),
    .Y(_1821_));
 sky130_fd_sc_hd__xor2_1 _6166_ (.A(_2822_),
    .B(_1821_),
    .X(_2711_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_2717_),
    .B(_2852_),
    .Y(_1822_));
 sky130_fd_sc_hd__o21ai_1 _6168_ (.A1(_2715_),
    .A2(_2852_),
    .B1(_1822_),
    .Y(_2137_));
 sky130_fd_sc_hd__o211ai_1 _6169_ (.A1(_2756_),
    .A2(_1817_),
    .B1(_0782_),
    .C1(net23),
    .Y(_1823_));
 sky130_fd_sc_hd__o21ai_0 _6170_ (.A1(net23),
    .A2(_0782_),
    .B1(_1823_),
    .Y(_2740_));
 sky130_fd_sc_hd__inv_1 _6171_ (.A(_0571_),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _6172_ (.A(_0592_),
    .B(_0594_),
    .Y(_1824_));
 sky130_fd_sc_hd__nor2_1 _6173_ (.A(_2640_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__nor2_1 _6174_ (.A(_0595_),
    .B(_1825_),
    .Y(_2834_));
 sky130_fd_sc_hd__xor2_1 _6175_ (.A(_2134_),
    .B(_2644_),
    .X(_2838_));
 sky130_fd_sc_hd__nor2_1 _6176_ (.A(_3057_),
    .B(_1750_),
    .Y(_1826_));
 sky130_fd_sc_hd__xor2_1 _6177_ (.A(_3034_),
    .B(_1826_),
    .X(_2900_));
 sky130_fd_sc_hd__o21ai_0 _6178_ (.A1(_2996_),
    .A2(_1749_),
    .B1(_0972_),
    .Y(_1827_));
 sky130_fd_sc_hd__xnor2_1 _6179_ (.A(_2992_),
    .B(_1827_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand2_1 _6180_ (.A(net26),
    .B(_1101_),
    .Y(_1828_));
 sky130_fd_sc_hd__xnor2_1 _6181_ (.A(_2996_),
    .B(_1828_),
    .Y(_2911_));
 sky130_fd_sc_hd__nor2_1 _6182_ (.A(_2920_),
    .B(_3057_),
    .Y(_1829_));
 sky130_fd_sc_hd__xor2_1 _6183_ (.A(_3000_),
    .B(_1829_),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(_2921_),
    .B(net26),
    .Y(_1830_));
 sky130_fd_sc_hd__o21ai_1 _6185_ (.A1(_2919_),
    .A2(_3038_),
    .B1(_1830_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2_1 _6186_ (.A(_0843_),
    .B(_0845_),
    .Y(_1831_));
 sky130_fd_sc_hd__nor2_1 _6187_ (.A(_2832_),
    .B(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nor2_1 _6188_ (.A(_0846_),
    .B(_1832_),
    .Y(_3012_));
 sky130_fd_sc_hd__nand2_1 _6189_ (.A(_0828_),
    .B(_0830_),
    .Y(_1833_));
 sky130_fd_sc_hd__nor2_1 _6190_ (.A(_2836_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__nor2_1 _6191_ (.A(_0831_),
    .B(_1834_),
    .Y(_3016_));
 sky130_fd_sc_hd__xnor2_1 _6192_ (.A(_2840_),
    .B(_2143_),
    .Y(_3020_));
 sky130_fd_sc_hd__nor2_1 _6193_ (.A(_3159_),
    .B(_3209_),
    .Y(_1835_));
 sky130_fd_sc_hd__a21oi_1 _6194_ (.A1(_1235_),
    .A2(_1835_),
    .B1(_1049_),
    .Y(_1836_));
 sky130_fd_sc_hd__xor2_1 _6195_ (.A(_3205_),
    .B(_1836_),
    .X(_3093_));
 sky130_fd_sc_hd__nor2b_1 _6196_ (.A(_3209_),
    .B_N(_1746_),
    .Y(_1837_));
 sky130_fd_sc_hd__nor2_1 _6197_ (.A(_3235_),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__xor2_1 _6198_ (.A(_3159_),
    .B(_1838_),
    .X(_3097_));
 sky130_fd_sc_hd__nor2_1 _6199_ (.A(_1049_),
    .B(_1235_),
    .Y(_1839_));
 sky130_fd_sc_hd__xor2_1 _6200_ (.A(_3209_),
    .B(_1839_),
    .X(_3101_));
 sky130_fd_sc_hd__nor2_1 _6201_ (.A(_3110_),
    .B(_3235_),
    .Y(_1840_));
 sky130_fd_sc_hd__xor2_1 _6202_ (.A(_3163_),
    .B(_1840_),
    .X(_3105_));
 sky130_fd_sc_hd__nand2_1 _6203_ (.A(_3111_),
    .B(_3213_),
    .Y(_1841_));
 sky130_fd_sc_hd__o21ai_1 _6204_ (.A1(_3108_),
    .A2(_3213_),
    .B1(_1841_),
    .Y(_2157_));
 sky130_fd_sc_hd__xor2_1 _6205_ (.A(_3010_),
    .B(_0996_),
    .X(_3176_));
 sky130_fd_sc_hd__xor2_1 _6206_ (.A(_3014_),
    .B(_1010_),
    .X(_3180_));
 sky130_fd_sc_hd__xnor2_1 _6207_ (.A(_2152_),
    .B(_3022_),
    .Y(_3188_));
 sky130_fd_sc_hd__nor2b_1 _6208_ (.A(_3040_),
    .B_N(_3043_),
    .Y(_1842_));
 sky130_fd_sc_hd__inv_1 _6209_ (.A(_3040_),
    .Y(_1843_));
 sky130_fd_sc_hd__nor3_1 _6210_ (.A(_1843_),
    .B(_3042_),
    .C(_3045_),
    .Y(_1844_));
 sky130_fd_sc_hd__o21ai_0 _6211_ (.A1(_3067_),
    .A2(_1762_),
    .B1(_3065_),
    .Y(_1845_));
 sky130_fd_sc_hd__a21boi_0 _6212_ (.A1(_1031_),
    .A2(_1845_),
    .B1_N(_3062_),
    .Y(_1846_));
 sky130_fd_sc_hd__o21ai_0 _6213_ (.A1(_3061_),
    .A2(_1846_),
    .B1(_3059_),
    .Y(_1847_));
 sky130_fd_sc_hd__a21boi_0 _6214_ (.A1(_1030_),
    .A2(_1847_),
    .B1_N(_3055_),
    .Y(_1848_));
 sky130_fd_sc_hd__o21ai_0 _6215_ (.A1(_3054_),
    .A2(_1848_),
    .B1(_3052_),
    .Y(_1849_));
 sky130_fd_sc_hd__a21boi_0 _6216_ (.A1(_1029_),
    .A2(_1849_),
    .B1_N(_3049_),
    .Y(_1850_));
 sky130_fd_sc_hd__o21ai_0 _6217_ (.A1(_3048_),
    .A2(_1850_),
    .B1(_3046_),
    .Y(_1851_));
 sky130_fd_sc_hd__mux2i_1 _6218_ (.A0(_1842_),
    .A1(_1844_),
    .S(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__nor3_1 _6219_ (.A(_1843_),
    .B(_3043_),
    .C(_3042_),
    .Y(_1853_));
 sky130_fd_sc_hd__a221oi_1 _6220_ (.A1(_1843_),
    .A2(_3042_),
    .B1(_3045_),
    .B2(_1842_),
    .C1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(_1852_),
    .B(_1854_),
    .Y(_3214_));
 sky130_fd_sc_hd__nand2_1 _6222_ (.A(_1028_),
    .B(_1045_),
    .Y(_1855_));
 sky130_fd_sc_hd__nor2_1 _6223_ (.A(_3043_),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__nor2_1 _6224_ (.A(_1046_),
    .B(_1856_),
    .Y(_3217_));
 sky130_fd_sc_hd__nor2_1 _6225_ (.A(_3048_),
    .B(_1850_),
    .Y(_1857_));
 sky130_fd_sc_hd__xnor2_1 _6226_ (.A(_3046_),
    .B(_1857_),
    .Y(_3220_));
 sky130_fd_sc_hd__nand2_1 _6227_ (.A(_1029_),
    .B(_1043_),
    .Y(_1858_));
 sky130_fd_sc_hd__nor2_1 _6228_ (.A(_3049_),
    .B(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__nor2_1 _6229_ (.A(_1044_),
    .B(_1859_),
    .Y(_3223_));
 sky130_fd_sc_hd__nor2_1 _6230_ (.A(_3054_),
    .B(_1848_),
    .Y(_1860_));
 sky130_fd_sc_hd__xnor2_1 _6231_ (.A(_3052_),
    .B(_1860_),
    .Y(_3226_));
 sky130_fd_sc_hd__nand2_1 _6232_ (.A(_1030_),
    .B(_1041_),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _6233_ (.A(_3055_),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor2_1 _6234_ (.A(_1042_),
    .B(_1862_),
    .Y(_3229_));
 sky130_fd_sc_hd__nor2_1 _6235_ (.A(_3061_),
    .B(_1846_),
    .Y(_1863_));
 sky130_fd_sc_hd__xnor2_1 _6236_ (.A(_3059_),
    .B(_1863_),
    .Y(_3232_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_1031_),
    .B(_1039_),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _6238_ (.A(_3062_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_1 _6239_ (.A(_1040_),
    .B(_1865_),
    .Y(_3236_));
 sky130_fd_sc_hd__nand2_1 _6240_ (.A(_1032_),
    .B(_1037_),
    .Y(_1866_));
 sky130_fd_sc_hd__nor2_1 _6241_ (.A(_3068_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__nor2_1 _6242_ (.A(_1038_),
    .B(_1867_),
    .Y(_3242_));
 sky130_fd_sc_hd__nor2_1 _6243_ (.A(_3073_),
    .B(_1760_),
    .Y(_1868_));
 sky130_fd_sc_hd__xnor2_1 _6244_ (.A(_3071_),
    .B(_1868_),
    .Y(_3245_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(_1033_),
    .B(_1035_),
    .Y(_1869_));
 sky130_fd_sc_hd__nor2_1 _6246_ (.A(_3074_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__nor2_1 _6247_ (.A(_1036_),
    .B(_1870_),
    .Y(_3248_));
 sky130_fd_sc_hd__xor2_1 _6248_ (.A(_3077_),
    .B(_1758_),
    .X(_3251_));
 sky130_fd_sc_hd__a21oi_1 _6249_ (.A1(_1238_),
    .A2(_1746_),
    .B1(net11),
    .Y(_1871_));
 sky130_fd_sc_hd__xnor2_1 _6250_ (.A(_1234_),
    .B(_1871_),
    .Y(_3258_));
 sky130_fd_sc_hd__nor2_1 _6251_ (.A(_1186_),
    .B(_1771_),
    .Y(_1872_));
 sky130_fd_sc_hd__xor2_1 _6252_ (.A(_3361_),
    .B(_1872_),
    .X(_3266_));
 sky130_fd_sc_hd__xnor2_1 _6253_ (.A(_3095_),
    .B(_1062_),
    .Y(_3270_));
 sky130_fd_sc_hd__xnor2_1 _6254_ (.A(_3099_),
    .B(_1191_),
    .Y(_3274_));
 sky130_fd_sc_hd__xnor2_1 _6255_ (.A(_3103_),
    .B(_1060_),
    .Y(_3278_));
 sky130_fd_sc_hd__xor2_1 _6256_ (.A(_3107_),
    .B(_2158_),
    .X(_3282_));
 sky130_fd_sc_hd__or2_1 _6257_ (.A(_1231_),
    .B(_1232_),
    .X(_1873_));
 sky130_fd_sc_hd__a31oi_2 _6258_ (.A1(_1234_),
    .A2(_1238_),
    .A3(_1746_),
    .B1(net25),
    .Y(_1874_));
 sky130_fd_sc_hd__a21o_1 _6259_ (.A1(_1873_),
    .A2(_1874_),
    .B1(_1233_),
    .X(_3295_));
 sky130_fd_sc_hd__a21o_1 _6260_ (.A1(_1873_),
    .A2(_1874_),
    .B1(_1233_),
    .X(_3303_));
 sky130_fd_sc_hd__xnor2_1 _6261_ (.A(_1873_),
    .B(_1239_),
    .Y(_3307_));
 sky130_fd_sc_hd__a21o_1 _6262_ (.A1(_1873_),
    .A2(_1874_),
    .B1(_1233_),
    .X(_3299_));
 sky130_fd_sc_hd__or2_0 _6263_ (.A(_1233_),
    .B(_1240_),
    .X(_3317_));
 sky130_fd_sc_hd__xnor2_1 _6264_ (.A(_3182_),
    .B(_1143_),
    .Y(_3343_));
 sky130_fd_sc_hd__inv_1 _6265_ (.A(_3247_),
    .Y(_1875_));
 sky130_fd_sc_hd__inv_1 _6266_ (.A(_3253_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2_1 _6267_ (.A(net28),
    .B(_3080_),
    .Y(_1877_));
 sky130_fd_sc_hd__o31a_1 _6268_ (.A1(_3039_),
    .A2(_3080_),
    .A3(_1047_),
    .B1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__o21bai_1 _6269_ (.A1(_1876_),
    .A2(_1878_),
    .B1_N(_3252_),
    .Y(_1879_));
 sky130_fd_sc_hd__a21oi_1 _6270_ (.A1(_3250_),
    .A2(_1879_),
    .B1(_3249_),
    .Y(_1880_));
 sky130_fd_sc_hd__o21bai_1 _6271_ (.A1(_1875_),
    .A2(_1880_),
    .B1_N(_3246_),
    .Y(_1881_));
 sky130_fd_sc_hd__a21o_1 _6272_ (.A1(_3244_),
    .A2(_1881_),
    .B1(_3243_),
    .X(_1882_));
 sky130_fd_sc_hd__a21oi_1 _6273_ (.A1(_3241_),
    .A2(_1882_),
    .B1(_3240_),
    .Y(_1883_));
 sky130_fd_sc_hd__o21bai_1 _6274_ (.A1(_1169_),
    .A2(_1883_),
    .B1_N(_3237_),
    .Y(_1884_));
 sky130_fd_sc_hd__a21oi_1 _6275_ (.A1(_3234_),
    .A2(_1884_),
    .B1(_3233_),
    .Y(_1885_));
 sky130_fd_sc_hd__o21bai_1 _6276_ (.A1(_1168_),
    .A2(_1885_),
    .B1_N(_3230_),
    .Y(_1886_));
 sky130_fd_sc_hd__a21o_1 _6277_ (.A1(_3225_),
    .A2(_3227_),
    .B1(_3224_),
    .X(_1887_));
 sky130_fd_sc_hd__a31o_1 _6278_ (.A1(_3225_),
    .A2(_3228_),
    .A3(_1886_),
    .B1(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__a21o_1 _6279_ (.A1(_3222_),
    .A2(_1888_),
    .B1(_3221_),
    .X(_1889_));
 sky130_fd_sc_hd__a21oi_1 _6280_ (.A1(_3219_),
    .A2(_1889_),
    .B1(_3218_),
    .Y(_1890_));
 sky130_fd_sc_hd__xnor2_1 _6281_ (.A(_3216_),
    .B(_1890_),
    .Y(_3381_));
 sky130_fd_sc_hd__xnor2_1 _6282_ (.A(_3219_),
    .B(_1183_),
    .Y(_3384_));
 sky130_fd_sc_hd__xor2_1 _6283_ (.A(_3222_),
    .B(_1888_),
    .X(_3387_));
 sky130_fd_sc_hd__xnor2_1 _6284_ (.A(_3225_),
    .B(_1181_),
    .Y(_3390_));
 sky130_fd_sc_hd__xor2_1 _6285_ (.A(_3228_),
    .B(_1886_),
    .X(_3393_));
 sky130_fd_sc_hd__xnor2_1 _6286_ (.A(_3231_),
    .B(_1179_),
    .Y(_3396_));
 sky130_fd_sc_hd__xor2_1 _6287_ (.A(_3234_),
    .B(_1884_),
    .X(_3399_));
 sky130_fd_sc_hd__xnor2_1 _6288_ (.A(_3238_),
    .B(_1177_),
    .Y(_3402_));
 sky130_fd_sc_hd__xor2_1 _6289_ (.A(_3241_),
    .B(_1882_),
    .X(_3406_));
 sky130_fd_sc_hd__xnor2_1 _6290_ (.A(_3244_),
    .B(_1175_),
    .Y(_3409_));
 sky130_fd_sc_hd__xnor2_1 _6291_ (.A(_3247_),
    .B(_1880_),
    .Y(_3412_));
 sky130_fd_sc_hd__xnor2_1 _6292_ (.A(_3250_),
    .B(_1173_),
    .Y(_3415_));
 sky130_fd_sc_hd__xnor2_1 _6293_ (.A(_3253_),
    .B(_1878_),
    .Y(_3418_));
 sky130_fd_sc_hd__xor2_1 _6294_ (.A(net28),
    .B(_3256_),
    .X(_3421_));
 sky130_fd_sc_hd__nand2_1 _6295_ (.A(_1464_),
    .B(_1465_),
    .Y(_3425_));
 sky130_fd_sc_hd__nand2_1 _6296_ (.A(_1431_),
    .B(_1433_),
    .Y(_3434_));
 sky130_fd_sc_hd__nand2_1 _6297_ (.A(_1431_),
    .B(_1433_),
    .Y(_3437_));
 sky130_fd_sc_hd__xnor2_1 _6298_ (.A(_3276_),
    .B(_1201_),
    .Y(_3445_));
 sky130_fd_sc_hd__nor2_1 _6299_ (.A(_1319_),
    .B(_1357_),
    .Y(_1891_));
 sky130_fd_sc_hd__xor2_1 _6300_ (.A(_3641_),
    .B(_1891_),
    .X(_3449_));
 sky130_fd_sc_hd__xor2_1 _6301_ (.A(_2168_),
    .B(_3284_),
    .X(_3453_));
 sky130_fd_sc_hd__nand2_1 _6302_ (.A(_3620_),
    .B(_3489_),
    .Y(_1892_));
 sky130_fd_sc_hd__xnor2_1 _6303_ (.A(_1356_),
    .B(_1892_),
    .Y(_2188_));
 sky130_fd_sc_hd__mux2_1 _6304_ (.A0(_1773_),
    .A1(net8),
    .S(_1770_),
    .X(_3466_));
 sky130_fd_sc_hd__nand2_1 _6305_ (.A(_1431_),
    .B(_1433_),
    .Y(_3470_));
 sky130_fd_sc_hd__o21ai_2 _6306_ (.A1(_3443_),
    .A2(_3517_),
    .B1(_1431_),
    .Y(_3474_));
 sky130_fd_sc_hd__xnor2_1 _6307_ (.A(_3268_),
    .B(_1203_),
    .Y(_3478_));
 sky130_fd_sc_hd__xnor2_1 _6308_ (.A(_3272_),
    .B(_1335_),
    .Y(_3482_));
 sky130_fd_sc_hd__o211ai_1 _6309_ (.A1(_3394_),
    .A2(_1792_),
    .B1(_3389_),
    .C1(_3392_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand2_1 _6310_ (.A(_3389_),
    .B(_3391_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand3_1 _6311_ (.A(_1312_),
    .B(_1893_),
    .C(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__a21oi_1 _6312_ (.A1(_3386_),
    .A2(_1895_),
    .B1(_3385_),
    .Y(_1896_));
 sky130_fd_sc_hd__xnor2_1 _6313_ (.A(_3383_),
    .B(_1896_),
    .Y(_3490_));
 sky130_fd_sc_hd__xor2_1 _6314_ (.A(_3386_),
    .B(_1313_),
    .X(_3493_));
 sky130_fd_sc_hd__xnor2_1 _6315_ (.A(_3395_),
    .B(_1791_),
    .Y(_3502_));
 sky130_fd_sc_hd__xor2_1 _6316_ (.A(_3398_),
    .B(_1308_),
    .X(_3505_));
 sky130_fd_sc_hd__xnor2_1 _6317_ (.A(_3401_),
    .B(_1789_),
    .Y(_3508_));
 sky130_fd_sc_hd__nor2_1 _6318_ (.A(_3404_),
    .B(_1305_),
    .Y(_1897_));
 sky130_fd_sc_hd__nor2_1 _6319_ (.A(_1306_),
    .B(_1897_),
    .Y(_3511_));
 sky130_fd_sc_hd__xnor2_1 _6320_ (.A(_3408_),
    .B(_1787_),
    .Y(_3514_));
 sky130_fd_sc_hd__a211oi_1 _6321_ (.A1(_3414_),
    .A2(_1301_),
    .B1(_3413_),
    .C1(_3411_),
    .Y(_1898_));
 sky130_fd_sc_hd__nor2_1 _6322_ (.A(_1303_),
    .B(_1898_),
    .Y(_3518_));
 sky130_fd_sc_hd__xor2_2 _6323_ (.A(_2172_),
    .B(_3353_),
    .X(_3530_));
 sky130_fd_sc_hd__nand2_1 _6324_ (.A(_1464_),
    .B(_1465_),
    .Y(_3534_));
 sky130_fd_sc_hd__nand2_1 _6325_ (.A(_1431_),
    .B(_1433_),
    .Y(_3538_));
 sky130_fd_sc_hd__xnor2_1 _6326_ (.A(_2178_),
    .B(net133),
    .Y(_3542_));
 sky130_fd_sc_hd__xor2_2 _6327_ (.A(_3349_),
    .B(_1282_),
    .X(_3546_));
 sky130_fd_sc_hd__mux2_1 _6328_ (.A0(_1773_),
    .A1(net8),
    .S(_1770_),
    .X(_3550_));
 sky130_fd_sc_hd__and2_0 _6329_ (.A(_1398_),
    .B(_1503_),
    .X(_1899_));
 sky130_fd_sc_hd__xnor2_1 _6330_ (.A(_3736_),
    .B(_1899_),
    .Y(_3558_));
 sky130_fd_sc_hd__xnor2_2 _6331_ (.A(_3345_),
    .B(_1268_),
    .Y(_3562_));
 sky130_fd_sc_hd__nand2_1 _6332_ (.A(_1464_),
    .B(_1465_),
    .Y(_3566_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(_1431_),
    .B(_1433_),
    .Y(_3570_));
 sky130_fd_sc_hd__o21ai_0 _6334_ (.A1(_3736_),
    .A2(_1527_),
    .B1(_1555_),
    .Y(_1900_));
 sky130_fd_sc_hd__xor2_1 _6335_ (.A(_3740_),
    .B(_1900_),
    .X(_3574_));
 sky130_fd_sc_hd__nand2_1 _6336_ (.A(_3489_),
    .B(_1490_),
    .Y(_1901_));
 sky130_fd_sc_hd__xor2_1 _6337_ (.A(_3569_),
    .B(_1901_),
    .X(_3578_));
 sky130_fd_sc_hd__mux2_1 _6338_ (.A0(_1773_),
    .A1(net8),
    .S(_1770_),
    .X(_3582_));
 sky130_fd_sc_hd__nand2_1 _6339_ (.A(_1431_),
    .B(_1433_),
    .Y(_3586_));
 sky130_fd_sc_hd__o31ai_1 _6340_ (.A1(_3736_),
    .A2(_3740_),
    .A3(_1503_),
    .B1(_1555_),
    .Y(_1902_));
 sky130_fd_sc_hd__xor2_1 _6341_ (.A(_3743_),
    .B(_1902_),
    .X(_3590_));
 sky130_fd_sc_hd__xnor2_1 _6342_ (.A(_3585_),
    .B(_1475_),
    .Y(_3594_));
 sky130_fd_sc_hd__nor2_1 _6343_ (.A(_3600_),
    .B(_1397_),
    .Y(_1903_));
 sky130_fd_sc_hd__nor2_1 _6344_ (.A(_1507_),
    .B(_1903_),
    .Y(_3602_));
 sky130_fd_sc_hd__xnor2_1 _6345_ (.A(_3379_),
    .B(_1286_),
    .Y(_3610_));
 sky130_fd_sc_hd__xor2_2 _6346_ (.A(_3612_),
    .B(net222),
    .X(_3617_));
 sky130_fd_sc_hd__a21oi_1 _6347_ (.A1(_1505_),
    .A2(_3597_),
    .B1(_1507_),
    .Y(_3625_));
 sky130_fd_sc_hd__nor2_2 _6348_ (.A(_3674_),
    .B(_1397_),
    .Y(_1904_));
 sky130_fd_sc_hd__xnor2_1 _6349_ (.A(_1904_),
    .B(net190),
    .Y(_3690_));
 sky130_fd_sc_hd__nand2_2 _6350_ (.A(_1804_),
    .B(_1555_),
    .Y(_1905_));
 sky130_fd_sc_hd__xnor2_1 _6351_ (.A(_3653_),
    .B(_1905_),
    .Y(_3694_));
 sky130_fd_sc_hd__xnor2_2 _6352_ (.A(_3447_),
    .B(_1365_),
    .Y(_3698_));
 sky130_fd_sc_hd__xnor2_2 _6353_ (.A(_3484_),
    .B(_1347_),
    .Y(_3702_));
 sky130_fd_sc_hd__or4_4 _6354_ (.A(_3653_),
    .B(_3661_),
    .C(_3669_),
    .D(_1802_),
    .X(_3706_));
 sky130_fd_sc_hd__o21bai_1 _6355_ (.A1(_3708_),
    .A2(_1397_),
    .B1_N(_1806_),
    .Y(_3710_));
 sky130_fd_sc_hd__nand2_1 _6356_ (.A(_3705_),
    .B(_1807_),
    .Y(_3713_));
 sky130_fd_sc_hd__xnor2_1 _6357_ (.A(net116),
    .B(_1349_),
    .Y(_3717_));
 sky130_fd_sc_hd__and3_1 _6358_ (.A(_1398_),
    .B(net197),
    .C(_1568_),
    .X(_1906_));
 sky130_fd_sc_hd__a21o_1 _6359_ (.A1(_1906_),
    .A2(net201),
    .B1(_1806_),
    .X(_3721_));
 sky130_fd_sc_hd__o21bai_1 _6360_ (.A1(_1807_),
    .A2(_1808_),
    .B1_N(_1806_),
    .Y(_3725_));
 sky130_fd_sc_hd__a21o_1 _6361_ (.A1(_1906_),
    .A2(net201),
    .B1(_1806_),
    .X(_3729_));
 sky130_fd_sc_hd__o21bai_1 _6362_ (.A1(_1807_),
    .A2(_1808_),
    .B1_N(_1806_),
    .Y(_3733_));
 sky130_fd_sc_hd__a21o_1 _6363_ (.A1(_3707_),
    .A2(_1555_),
    .B1(_1806_),
    .X(_3744_));
 sky130_fd_sc_hd__inv_1 _6364_ (.A(_3526_),
    .Y(net94));
 sky130_fd_sc_hd__inv_1 _6365_ (.A(_3723_),
    .Y(_1907_));
 sky130_fd_sc_hd__inv_1 _6366_ (.A(_3712_),
    .Y(_1908_));
 sky130_fd_sc_hd__inv_1 _6367_ (.A(_3700_),
    .Y(_1909_));
 sky130_fd_sc_hd__inv_1 _6368_ (.A(_3696_),
    .Y(_1910_));
 sky130_fd_sc_hd__a21oi_2 _6369_ (.A1(_3692_),
    .A2(_2193_),
    .B1(_3691_),
    .Y(_1911_));
 sky130_fd_sc_hd__nor2_1 _6370_ (.A(_1911_),
    .B(_1910_),
    .Y(_1912_));
 sky130_fd_sc_hd__nor2_2 _6371_ (.A(_1912_),
    .B(_3695_),
    .Y(_1913_));
 sky130_fd_sc_hd__o21bai_1 _6372_ (.A1(_1909_),
    .A2(_1913_),
    .B1_N(_3699_),
    .Y(_1914_));
 sky130_fd_sc_hd__a21oi_2 _6373_ (.A1(_1914_),
    .A2(_3704_),
    .B1(_3703_),
    .Y(_1915_));
 sky130_fd_sc_hd__o21bai_1 _6374_ (.A1(_1915_),
    .A2(_1908_),
    .B1_N(_3711_),
    .Y(_1916_));
 sky130_fd_sc_hd__a21oi_2 _6375_ (.A1(_1916_),
    .A2(_3719_),
    .B1(_3718_),
    .Y(_1917_));
 sky130_fd_sc_hd__o21bai_1 _6376_ (.A1(_1917_),
    .A2(_1907_),
    .B1_N(_3722_),
    .Y(_1918_));
 sky130_fd_sc_hd__a21oi_2 _6377_ (.A1(_3727_),
    .A2(_1918_),
    .B1(_3726_),
    .Y(_1919_));
 sky130_fd_sc_hd__xnor2_2 _6378_ (.A(_3731_),
    .B(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__buf_2 _6379_ (.A(_3686_),
    .X(_1921_));
 sky130_fd_sc_hd__inv_1 _6380_ (.A(_3719_),
    .Y(_1922_));
 sky130_fd_sc_hd__inv_1 _6381_ (.A(_3704_),
    .Y(_1923_));
 sky130_fd_sc_hd__a21o_1 _6382_ (.A1(_3677_),
    .A2(_2191_),
    .B1(_3676_),
    .X(_1924_));
 sky130_fd_sc_hd__a21oi_2 _6383_ (.A1(_1924_),
    .A2(_3692_),
    .B1(_3691_),
    .Y(_1925_));
 sky130_fd_sc_hd__o21bai_1 _6384_ (.A1(_1925_),
    .A2(_1910_),
    .B1_N(_3695_),
    .Y(_1926_));
 sky130_fd_sc_hd__a21oi_2 _6385_ (.A1(_1926_),
    .A2(_3700_),
    .B1(_3699_),
    .Y(_1927_));
 sky130_fd_sc_hd__o21bai_1 _6386_ (.A1(_1923_),
    .A2(_1927_),
    .B1_N(_3703_),
    .Y(_1928_));
 sky130_fd_sc_hd__a21oi_2 _6387_ (.A1(_3712_),
    .A2(_1928_),
    .B1(_3711_),
    .Y(_1929_));
 sky130_fd_sc_hd__o21bai_1 _6388_ (.A1(_1922_),
    .A2(_1929_),
    .B1_N(_3718_),
    .Y(_1930_));
 sky130_fd_sc_hd__a21oi_4 _6389_ (.A1(_3723_),
    .A2(_1930_),
    .B1(_3722_),
    .Y(_1931_));
 sky130_fd_sc_hd__xnor2_2 _6390_ (.A(_3727_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__xnor2_2 _6391_ (.A(net208),
    .B(_3723_),
    .Y(_1933_));
 sky130_fd_sc_hd__xnor2_2 _6392_ (.A(net221),
    .B(_3719_),
    .Y(_1934_));
 sky130_fd_sc_hd__xnor2_2 _6393_ (.A(_1915_),
    .B(_3712_),
    .Y(_1935_));
 sky130_fd_sc_hd__xnor2_4 _6394_ (.A(_1923_),
    .B(net233),
    .Y(_1936_));
 sky130_fd_sc_hd__xnor2_2 _6395_ (.A(_3700_),
    .B(_1913_),
    .Y(_1937_));
 sky130_fd_sc_hd__xnor2_4 _6396_ (.A(net228),
    .B(net209),
    .Y(_1938_));
 sky130_fd_sc_hd__nor2_2 _6397_ (.A(_1937_),
    .B(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__xnor2_4 _6398_ (.A(_3692_),
    .B(net129),
    .Y(_1940_));
 sky130_fd_sc_hd__nand4_1 _6399_ (.A(_3681_),
    .B(_1936_),
    .C(_1939_),
    .D(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__or3_4 _6400_ (.A(_1941_),
    .B(net210),
    .C(_1934_),
    .X(_1942_));
 sky130_fd_sc_hd__or3_4 _6401_ (.A(_1932_),
    .B(_1942_),
    .C(_1933_),
    .X(_1943_));
 sky130_fd_sc_hd__nand2_4 _6402_ (.A(_1943_),
    .B(_1921_),
    .Y(_1944_));
 sky130_fd_sc_hd__xnor2_2 _6403_ (.A(_1920_),
    .B(_1944_),
    .Y(net79));
 sky130_fd_sc_hd__inv_1 _6404_ (.A(_3727_),
    .Y(_1945_));
 sky130_fd_sc_hd__o21bai_1 _6405_ (.A1(_1945_),
    .A2(_1931_),
    .B1_N(_3726_),
    .Y(_1946_));
 sky130_fd_sc_hd__a21oi_2 _6406_ (.A1(_3731_),
    .A2(_1946_),
    .B1(_3730_),
    .Y(_1947_));
 sky130_fd_sc_hd__xnor2_2 _6407_ (.A(_3735_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nor2_1 _6408_ (.A(net78),
    .B(_2194_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand3_2 _6409_ (.A(_1939_),
    .B(_1940_),
    .C(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__or3b_4 _6410_ (.A(_1950_),
    .B(_1935_),
    .C_N(_1936_),
    .X(_1951_));
 sky130_fd_sc_hd__or3_4 _6411_ (.A(_1951_),
    .B(_1934_),
    .C(_1933_),
    .X(_1952_));
 sky130_fd_sc_hd__or3_4 _6412_ (.A(_1920_),
    .B(_1952_),
    .C(_1932_),
    .X(_1953_));
 sky130_fd_sc_hd__nand2_2 _6413_ (.A(_1953_),
    .B(_1921_),
    .Y(_1954_));
 sky130_fd_sc_hd__xnor2_1 _6414_ (.A(_1948_),
    .B(_1954_),
    .Y(net80));
 sky130_fd_sc_hd__inv_1 _6415_ (.A(_3731_),
    .Y(_1955_));
 sky130_fd_sc_hd__o21bai_1 _6416_ (.A1(_1919_),
    .A2(_1955_),
    .B1_N(_3730_),
    .Y(_1956_));
 sky130_fd_sc_hd__a21oi_2 _6417_ (.A1(_1956_),
    .A2(_3735_),
    .B1(_3734_),
    .Y(_1957_));
 sky130_fd_sc_hd__xnor2_2 _6418_ (.A(_3738_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__or3_4 _6419_ (.A(_1920_),
    .B(_1943_),
    .C(_1948_),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_4 _6420_ (.A(_1959_),
    .B(_1921_),
    .Y(_1960_));
 sky130_fd_sc_hd__xnor2_2 _6421_ (.A(_1958_),
    .B(_1960_),
    .Y(net81));
 sky130_fd_sc_hd__inv_1 _6422_ (.A(_3735_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21bai_1 _6423_ (.A1(_1961_),
    .A2(_1947_),
    .B1_N(_3734_),
    .Y(_1962_));
 sky130_fd_sc_hd__a21oi_1 _6424_ (.A1(_3738_),
    .A2(_1962_),
    .B1(_3737_),
    .Y(_1963_));
 sky130_fd_sc_hd__xnor2_2 _6425_ (.A(_3742_),
    .B(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__o31ai_4 _6426_ (.A1(_1948_),
    .A2(_1958_),
    .A3(_1953_),
    .B1(_3686_),
    .Y(_1965_));
 sky130_fd_sc_hd__xnor2_2 _6427_ (.A(_1964_),
    .B(net119),
    .Y(net82));
 sky130_fd_sc_hd__inv_1 _6428_ (.A(_3738_),
    .Y(_1966_));
 sky130_fd_sc_hd__o21bai_1 _6429_ (.A1(_1957_),
    .A2(_1966_),
    .B1_N(_3737_),
    .Y(_1967_));
 sky130_fd_sc_hd__a21oi_1 _6430_ (.A1(_1967_),
    .A2(_3742_),
    .B1(_3741_),
    .Y(_1968_));
 sky130_fd_sc_hd__xnor2_1 _6431_ (.A(_1968_),
    .B(_3746_),
    .Y(_1969_));
 sky130_fd_sc_hd__o31ai_4 _6432_ (.A1(_1958_),
    .A2(_1964_),
    .A3(_1959_),
    .B1(_3686_),
    .Y(_1970_));
 sky130_fd_sc_hd__xnor2_1 _6433_ (.A(net196),
    .B(_1970_),
    .Y(net83));
 sky130_fd_sc_hd__a31oi_2 _6434_ (.A1(_3588_),
    .A2(_1482_),
    .A3(_1484_),
    .B1(_3587_),
    .Y(_1971_));
 sky130_fd_sc_hd__o21ai_1 _6435_ (.A1(_1964_),
    .A2(_1969_),
    .B1(_3686_),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2_1 _6436_ (.A(_1965_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__inv_1 _6437_ (.A(_3742_),
    .Y(_1974_));
 sky130_fd_sc_hd__o21bai_1 _6438_ (.A1(_1974_),
    .A2(_1963_),
    .B1_N(_3741_),
    .Y(_1975_));
 sky130_fd_sc_hd__a21oi_1 _6439_ (.A1(_3746_),
    .A2(_1975_),
    .B1(_3745_),
    .Y(_1976_));
 sky130_fd_sc_hd__xor2_1 _6440_ (.A(_1976_),
    .B(_1973_),
    .X(_1977_));
 sky130_fd_sc_hd__xnor3_1 _6441_ (.A(_1480_),
    .B(_1971_),
    .C(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__nor2_1 _6442_ (.A(_3714_),
    .B(_1397_),
    .Y(_1979_));
 sky130_fd_sc_hd__a31oi_2 _6443_ (.A1(_1397_),
    .A2(net198),
    .A3(_1568_),
    .B1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__xnor2_1 _6444_ (.A(_1978_),
    .B(_1980_),
    .Y(net84));
 sky130_fd_sc_hd__nand2_2 _6445_ (.A(_1921_),
    .B(_3682_),
    .Y(_1981_));
 sky130_fd_sc_hd__o21ai_2 _6446_ (.A1(_3679_),
    .A2(_1921_),
    .B1(_1981_),
    .Y(net85));
 sky130_fd_sc_hd__nor2b_2 _6447_ (.A(_3681_),
    .B_N(_3686_),
    .Y(_1982_));
 sky130_fd_sc_hd__xnor2_1 _6448_ (.A(_1982_),
    .B(net236),
    .Y(net86));
 sky130_fd_sc_hd__nand2_1 _6449_ (.A(_1940_),
    .B(_1949_),
    .Y(_1983_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_1921_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__xnor2_1 _6451_ (.A(_1984_),
    .B(_1938_),
    .Y(net87));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(_3681_),
    .B(net235),
    .Y(_1985_));
 sky130_fd_sc_hd__o21ai_2 _6453_ (.A1(_1985_),
    .A2(_1938_),
    .B1(_3686_),
    .Y(_1986_));
 sky130_fd_sc_hd__xnor2_1 _6454_ (.A(_1986_),
    .B(_1937_),
    .Y(net88));
 sky130_fd_sc_hd__nand2_1 _6455_ (.A(_1950_),
    .B(_3686_),
    .Y(_1987_));
 sky130_fd_sc_hd__xor2_1 _6456_ (.A(_1987_),
    .B(net229),
    .X(net89));
 sky130_fd_sc_hd__nand2_1 _6457_ (.A(_1921_),
    .B(_1941_),
    .Y(_1988_));
 sky130_fd_sc_hd__xnor2_2 _6458_ (.A(_1988_),
    .B(net210),
    .Y(net90));
 sky130_fd_sc_hd__nand2_2 _6459_ (.A(_1951_),
    .B(_1921_),
    .Y(_1989_));
 sky130_fd_sc_hd__xnor2_1 _6460_ (.A(_1934_),
    .B(_1989_),
    .Y(net91));
 sky130_fd_sc_hd__nand2_2 _6461_ (.A(_1942_),
    .B(_1921_),
    .Y(_1990_));
 sky130_fd_sc_hd__xnor2_1 _6462_ (.A(_1933_),
    .B(_1990_),
    .Y(net92));
 sky130_fd_sc_hd__nand2_2 _6463_ (.A(_1952_),
    .B(_1921_),
    .Y(_1991_));
 sky130_fd_sc_hd__xnor2_1 _6464_ (.A(_1932_),
    .B(_1991_),
    .Y(net93));
 sky130_fd_sc_hd__nor2b_1 _6465_ (.A(_2183_),
    .B_N(_3544_),
    .Y(_1992_));
 sky130_fd_sc_hd__o21ai_1 _6466_ (.A1(_3543_),
    .A2(_1992_),
    .B1(_3560_),
    .Y(_1993_));
 sky130_fd_sc_hd__nand2b_1 _6467_ (.A_N(_3559_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__a21o_1 _6468_ (.A1(_3576_),
    .A2(_1994_),
    .B1(_3575_),
    .X(_1995_));
 sky130_fd_sc_hd__a21o_1 _6469_ (.A1(_3592_),
    .A2(_1995_),
    .B1(_3591_),
    .X(_1996_));
 sky130_fd_sc_hd__a21o_1 _6470_ (.A1(_3604_),
    .A2(_1996_),
    .B1(_3603_),
    .X(_1997_));
 sky130_fd_sc_hd__a21o_1 _6471_ (.A1(_1997_),
    .A2(_3619_),
    .B1(_3618_),
    .X(_1998_));
 sky130_fd_sc_hd__a21o_1 _6472_ (.A1(_3627_),
    .A2(_1998_),
    .B1(_3626_),
    .X(_1999_));
 sky130_fd_sc_hd__a21oi_2 _6473_ (.A1(_1999_),
    .A2(_3631_),
    .B1(_3630_),
    .Y(_2000_));
 sky130_fd_sc_hd__xnor2_4 _6474_ (.A(_3639_),
    .B(net120),
    .Y(_2001_));
 sky130_fd_sc_hd__nor2_1 _6475_ (.A(_3684_),
    .B(_3685_),
    .Y(_2002_));
 sky130_fd_sc_hd__clkbuf_2 _6476_ (.A(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__nor2b_1 _6477_ (.A(_2181_),
    .B_N(_3525_),
    .Y(_2004_));
 sky130_fd_sc_hd__o21ai_1 _6478_ (.A1(_3524_),
    .A2(_2004_),
    .B1(_3544_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2b_1 _6479_ (.A_N(_3543_),
    .B(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__a21o_1 _6480_ (.A1(_3560_),
    .A2(_2006_),
    .B1(_3559_),
    .X(_2007_));
 sky130_fd_sc_hd__a21oi_2 _6481_ (.A1(_3576_),
    .A2(_2007_),
    .B1(_3575_),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2b_1 _6482_ (.A(_2008_),
    .B_N(_3592_),
    .Y(_2009_));
 sky130_fd_sc_hd__o21ai_1 _6483_ (.A1(_3591_),
    .A2(_2009_),
    .B1(_3604_),
    .Y(_2010_));
 sky130_fd_sc_hd__nand2b_1 _6484_ (.A_N(_3603_),
    .B(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__a21o_1 _6485_ (.A1(_3619_),
    .A2(_2011_),
    .B1(_3618_),
    .X(_2012_));
 sky130_fd_sc_hd__a21o_1 _6486_ (.A1(_2012_),
    .A2(_3627_),
    .B1(_3626_),
    .X(_2013_));
 sky130_fd_sc_hd__xor2_2 _6487_ (.A(_3631_),
    .B(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__xor2_1 _6488_ (.A(_3627_),
    .B(_1998_),
    .X(_2015_));
 sky130_fd_sc_hd__xor2_1 _6489_ (.A(_3619_),
    .B(_2011_),
    .X(_2016_));
 sky130_fd_sc_hd__xor2_1 _6490_ (.A(_3604_),
    .B(_1996_),
    .X(_2017_));
 sky130_fd_sc_hd__xnor2_2 _6491_ (.A(_3592_),
    .B(_2008_),
    .Y(_2018_));
 sky130_fd_sc_hd__xor2_4 _6492_ (.A(_3576_),
    .B(net142),
    .X(_2019_));
 sky130_fd_sc_hd__xor2_4 _6493_ (.A(net152),
    .B(net173),
    .X(_2020_));
 sky130_fd_sc_hd__xor2_4 _6494_ (.A(net144),
    .B(net240),
    .X(_2021_));
 sky130_fd_sc_hd__nand2_1 _6495_ (.A(_2021_),
    .B(_3527_),
    .Y(_2022_));
 sky130_fd_sc_hd__or4_1 _6496_ (.A(_2022_),
    .B(_2019_),
    .C(_2020_),
    .D(_2018_),
    .X(_2023_));
 sky130_fd_sc_hd__or3_1 _6497_ (.A(_2016_),
    .B(_2017_),
    .C(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__or3_4 _6498_ (.A(_2024_),
    .B(_2015_),
    .C(_2014_),
    .X(_2025_));
 sky130_fd_sc_hd__nand2_2 _6499_ (.A(_2003_),
    .B(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__xnor2_1 _6500_ (.A(_2001_),
    .B(_2026_),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _6501_ (.A(_3639_),
    .Y(_2027_));
 sky130_fd_sc_hd__a21oi_2 _6502_ (.A1(_2013_),
    .A2(_3631_),
    .B1(_3630_),
    .Y(_2028_));
 sky130_fd_sc_hd__o21bai_4 _6503_ (.A1(_2028_),
    .A2(_2027_),
    .B1_N(_3638_),
    .Y(_2029_));
 sky130_fd_sc_hd__xor2_4 _6504_ (.A(_2029_),
    .B(_3647_),
    .X(_2030_));
 sky130_fd_sc_hd__nor2_1 _6505_ (.A(_2019_),
    .B(_2020_),
    .Y(_2031_));
 sky130_fd_sc_hd__nand4_1 _6506_ (.A(_2031_),
    .B(_3526_),
    .C(_2184_),
    .D(_2021_),
    .Y(_2032_));
 sky130_fd_sc_hd__or3_1 _6507_ (.A(_2017_),
    .B(_2018_),
    .C(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__or3_4 _6508_ (.A(_2015_),
    .B(_2016_),
    .C(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__o31ai_4 _6509_ (.A1(_2001_),
    .A2(_2014_),
    .A3(_2034_),
    .B1(_2003_),
    .Y(_2035_));
 sky130_fd_sc_hd__xnor2_2 _6510_ (.A(_2035_),
    .B(_2030_),
    .Y(net96));
 sky130_fd_sc_hd__o21bai_1 _6511_ (.A1(_2027_),
    .A2(_2000_),
    .B1_N(_3638_),
    .Y(_2036_));
 sky130_fd_sc_hd__a21o_1 _6512_ (.A1(_2036_),
    .A2(_3647_),
    .B1(_3646_),
    .X(_2037_));
 sky130_fd_sc_hd__xor2_2 _6513_ (.A(_3655_),
    .B(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__o31ai_2 _6514_ (.A1(_2001_),
    .A2(_2025_),
    .A3(_2030_),
    .B1(_2003_),
    .Y(_2039_));
 sky130_fd_sc_hd__xnor2_1 _6515_ (.A(_2038_),
    .B(_2039_),
    .Y(net97));
 sky130_fd_sc_hd__a21o_1 _6516_ (.A1(_3647_),
    .A2(_2029_),
    .B1(_3646_),
    .X(_2040_));
 sky130_fd_sc_hd__a21oi_2 _6517_ (.A1(_2040_),
    .A2(_3655_),
    .B1(_3654_),
    .Y(_2041_));
 sky130_fd_sc_hd__xnor2_2 _6518_ (.A(_3663_),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__or4_4 _6519_ (.A(_2001_),
    .B(_2014_),
    .C(_2034_),
    .D(_2038_),
    .X(_2043_));
 sky130_fd_sc_hd__o21ai_4 _6520_ (.A1(_2043_),
    .A2(_2030_),
    .B1(_2002_),
    .Y(_2044_));
 sky130_fd_sc_hd__xnor2_1 _6521_ (.A(_2042_),
    .B(_2044_),
    .Y(net98));
 sky130_fd_sc_hd__inv_1 _6522_ (.A(_3663_),
    .Y(_2045_));
 sky130_fd_sc_hd__a21oi_1 _6523_ (.A1(_3655_),
    .A2(_2037_),
    .B1(_3654_),
    .Y(_2046_));
 sky130_fd_sc_hd__nor2_1 _6524_ (.A(_2045_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__nor2_1 _6525_ (.A(_3662_),
    .B(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__xnor2_1 _6526_ (.A(_3671_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__or4_1 _6527_ (.A(_2001_),
    .B(_2025_),
    .C(_2030_),
    .D(_2038_),
    .X(_2050_));
 sky130_fd_sc_hd__o21ai_2 _6528_ (.A1(_2042_),
    .A2(_2050_),
    .B1(_2003_),
    .Y(_2051_));
 sky130_fd_sc_hd__xnor2_1 _6529_ (.A(_2051_),
    .B(_2049_),
    .Y(net99));
 sky130_fd_sc_hd__o21bai_1 _6530_ (.A1(_2045_),
    .A2(_2041_),
    .B1_N(_3662_),
    .Y(_2052_));
 sky130_fd_sc_hd__a21oi_1 _6531_ (.A1(_3671_),
    .A2(_2052_),
    .B1(_3670_),
    .Y(_2053_));
 sky130_fd_sc_hd__o21ai_1 _6532_ (.A1(_2042_),
    .A2(_2049_),
    .B1(_2002_),
    .Y(_2054_));
 sky130_fd_sc_hd__nand2_2 _6533_ (.A(_2044_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__xnor2_2 _6534_ (.A(_2055_),
    .B(_2053_),
    .Y(_2056_));
 sky130_fd_sc_hd__nor2_1 _6535_ (.A(_3587_),
    .B(_1398_),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _6536_ (.A(_1480_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__nor3_1 _6537_ (.A(_3571_),
    .B(_1447_),
    .C(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__nand2_1 _6538_ (.A(_3588_),
    .B(_1396_),
    .Y(_2060_));
 sky130_fd_sc_hd__nor4b_1 _6539_ (.A(_1480_),
    .B(_1483_),
    .C(_2060_),
    .D_N(_1482_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _6540_ (.A(_3587_),
    .B(_1396_),
    .Y(_2062_));
 sky130_fd_sc_hd__nor2_1 _6541_ (.A(_3588_),
    .B(_3587_),
    .Y(_2063_));
 sky130_fd_sc_hd__nand3_1 _6542_ (.A(_1396_),
    .B(_1480_),
    .C(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_3614_),
    .B(_1398_),
    .Y(_2065_));
 sky130_fd_sc_hd__o211ai_1 _6544_ (.A1(_1480_),
    .A2(_2062_),
    .B1(_2064_),
    .C1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__nor3_1 _6545_ (.A(_2059_),
    .B(_2061_),
    .C(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__xnor3_1 _6546_ (.A(_3705_),
    .B(_2067_),
    .C(_2056_),
    .X(net100));
 sky130_fd_sc_hd__nand2b_1 _6547_ (.A_N(_3685_),
    .B(net68),
    .Y(_2068_));
 sky130_fd_sc_hd__nor2_2 _6548_ (.A(_3528_),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__a21oi_1 _6549_ (.A1(_2184_),
    .A2(_2068_),
    .B1(_2069_),
    .Y(net101));
 sky130_fd_sc_hd__nor2_1 _6550_ (.A(_3527_),
    .B(_2068_),
    .Y(_2070_));
 sky130_fd_sc_hd__xnor2_1 _6551_ (.A(net242),
    .B(_2070_),
    .Y(net102));
 sky130_fd_sc_hd__a31oi_1 _6552_ (.A1(net241),
    .A2(_3526_),
    .A3(_2184_),
    .B1(_2068_),
    .Y(_2071_));
 sky130_fd_sc_hd__xor2_1 _6553_ (.A(_2020_),
    .B(_2071_),
    .X(net103));
 sky130_fd_sc_hd__o21ai_2 _6554_ (.A1(_2022_),
    .A2(_2020_),
    .B1(_2003_),
    .Y(_2072_));
 sky130_fd_sc_hd__xnor2_1 _6555_ (.A(_2019_),
    .B(_2072_),
    .Y(net104));
 sky130_fd_sc_hd__nand2_1 _6556_ (.A(_2003_),
    .B(_2032_),
    .Y(_2073_));
 sky130_fd_sc_hd__xnor2_2 _6557_ (.A(net215),
    .B(_2073_),
    .Y(net105));
 sky130_fd_sc_hd__nand2_1 _6558_ (.A(_2003_),
    .B(_2023_),
    .Y(_2074_));
 sky130_fd_sc_hd__xnor2_1 _6559_ (.A(_2017_),
    .B(_2074_),
    .Y(net106));
 sky130_fd_sc_hd__nand2_2 _6560_ (.A(_2003_),
    .B(_2033_),
    .Y(_2075_));
 sky130_fd_sc_hd__xnor2_2 _6561_ (.A(_2016_),
    .B(_2075_),
    .Y(net107));
 sky130_fd_sc_hd__nand2_2 _6562_ (.A(_2003_),
    .B(_2024_),
    .Y(_2076_));
 sky130_fd_sc_hd__xnor2_2 _6563_ (.A(_2015_),
    .B(_2076_),
    .Y(net108));
 sky130_fd_sc_hd__nand2_2 _6564_ (.A(_2003_),
    .B(_2034_),
    .Y(_2077_));
 sky130_fd_sc_hd__xnor2_1 _6565_ (.A(_2014_),
    .B(_2077_),
    .Y(net109));
 sky130_fd_sc_hd__fa_4 _6566_ (.A(_2078_),
    .B(net53),
    .CIN(_2079_),
    .COUT(_2080_),
    .SUM(_2081_));
 sky130_fd_sc_hd__fa_4 _6567_ (.A(_2078_),
    .B(_2082_),
    .CIN(_2083_),
    .COUT(_2084_),
    .SUM(_2085_));
 sky130_fd_sc_hd__fa_2 _6568_ (.A(net37),
    .B(_2082_),
    .CIN(_2086_),
    .COUT(_2087_),
    .SUM(_2088_));
 sky130_fd_sc_hd__fa_4 _6569_ (.A(_2090_),
    .B(_2089_),
    .CIN(_2091_),
    .COUT(_2092_),
    .SUM(_2093_));
 sky130_fd_sc_hd__fa_2 _6570_ (.A(_2094_),
    .B(_2095_),
    .CIN(_2096_),
    .COUT(_2097_),
    .SUM(_2098_));
 sky130_fd_sc_hd__fa_1 _6571_ (.A(_2099_),
    .B(_2100_),
    .CIN(_2101_),
    .COUT(_2102_),
    .SUM(_2103_));
 sky130_fd_sc_hd__fa_1 _6572_ (.A(_2106_),
    .B(_2107_),
    .CIN(net5),
    .COUT(_2108_),
    .SUM(_2109_));
 sky130_fd_sc_hd__fa_1 _6573_ (.A(_2112_),
    .B(_2098_),
    .CIN(_2113_),
    .COUT(_2114_),
    .SUM(_2115_));
 sky130_fd_sc_hd__fa_1 _6574_ (.A(_2116_),
    .B(_2117_),
    .CIN(_2118_),
    .COUT(_2119_),
    .SUM(_2120_));
 sky130_fd_sc_hd__fa_1 _6575_ (.A(_2122_),
    .B(_2123_),
    .CIN(_2124_),
    .COUT(_2125_),
    .SUM(_2126_));
 sky130_fd_sc_hd__fa_1 _6576_ (.A(_2127_),
    .B(_2115_),
    .CIN(_2128_),
    .COUT(_2129_),
    .SUM(_2130_));
 sky130_fd_sc_hd__fa_1 _6577_ (.A(_2131_),
    .B(_2132_),
    .CIN(_2133_),
    .COUT(_2134_),
    .SUM(_2135_));
 sky130_fd_sc_hd__fa_1 _6578_ (.A(_2136_),
    .B(_2130_),
    .CIN(_2137_),
    .COUT(_2138_),
    .SUM(_2139_));
 sky130_fd_sc_hd__fa_1 _6579_ (.A(_2140_),
    .B(_2141_),
    .CIN(_2142_),
    .COUT(_2143_),
    .SUM(_2144_));
 sky130_fd_sc_hd__fa_4 _6580_ (.A(_2146_),
    .B(_2139_),
    .CIN(_2147_),
    .COUT(_2148_),
    .SUM(_2149_));
 sky130_fd_sc_hd__fa_1 _6581_ (.A(_2144_),
    .B(_2150_),
    .CIN(_2151_),
    .COUT(_2152_),
    .SUM(_2153_));
 sky130_fd_sc_hd__fa_1 _6582_ (.A(_2156_),
    .B(_2149_),
    .CIN(_2157_),
    .COUT(_2158_),
    .SUM(_2159_));
 sky130_fd_sc_hd__fa_1 _6583_ (.A(_2160_),
    .B(_2161_),
    .CIN(_2162_),
    .COUT(_2163_),
    .SUM(_2164_));
 sky130_fd_sc_hd__fa_2 _6584_ (.A(_2166_),
    .B(_2167_),
    .CIN(_2159_),
    .COUT(_2168_),
    .SUM(_2169_));
 sky130_fd_sc_hd__fa_2 _6585_ (.A(_2164_),
    .B(_2170_),
    .CIN(_2171_),
    .COUT(_2172_),
    .SUM(_2173_));
 sky130_fd_sc_hd__fa_2 _6586_ (.A(_2175_),
    .B(_2176_),
    .CIN(_2177_),
    .COUT(_2178_),
    .SUM(_2179_));
 sky130_fd_sc_hd__fa_2 _6587_ (.A(_2179_),
    .B(_2181_),
    .CIN(_2182_),
    .COUT(_2183_),
    .SUM(_2184_));
 sky130_fd_sc_hd__fa_2 _6588_ (.A(_2169_),
    .B(_2187_),
    .CIN(_2188_),
    .COUT(_2189_),
    .SUM(_2190_));
 sky130_fd_sc_hd__fa_2 _6589_ (.A(_2192_),
    .B(_2191_),
    .CIN(_2190_),
    .COUT(_2193_),
    .SUM(_2194_));
 sky130_fd_sc_hd__ha_1 _6590_ (.A(_2195_),
    .B(net46),
    .COUT(_2079_),
    .SUM(_2196_));
 sky130_fd_sc_hd__ha_1 _6591_ (.A(net30),
    .B(_2197_),
    .COUT(_2086_),
    .SUM(_2198_));
 sky130_fd_sc_hd__ha_1 _6592_ (.A(net30),
    .B(net46),
    .COUT(_2199_),
    .SUM(_2200_));
 sky130_fd_sc_hd__ha_1 _6593_ (.A(_2078_),
    .B(net53),
    .COUT(_2202_),
    .SUM(_2201_));
 sky130_fd_sc_hd__ha_1 _6594_ (.A(net37),
    .B(_2082_),
    .COUT(_2203_),
    .SUM(_2204_));
 sky130_fd_sc_hd__ha_1 _6595_ (.A(net37),
    .B(net53),
    .COUT(_2205_),
    .SUM(_2206_));
 sky130_fd_sc_hd__ha_1 _6596_ (.A(_2207_),
    .B(_2196_),
    .COUT(_2104_),
    .SUM(_2208_));
 sky130_fd_sc_hd__ha_2 _6597_ (.A(_2209_),
    .B(net55),
    .COUT(_2210_),
    .SUM(_2211_));
 sky130_fd_sc_hd__ha_2 _6598_ (.A(net39),
    .B(_2212_),
    .COUT(_2213_),
    .SUM(_2214_));
 sky130_fd_sc_hd__ha_1 _6599_ (.A(net39),
    .B(net55),
    .COUT(_2215_),
    .SUM(_2216_));
 sky130_fd_sc_hd__ha_1 _6600_ (.A(_2217_),
    .B(net54),
    .COUT(_2218_),
    .SUM(_2219_));
 sky130_fd_sc_hd__ha_2 _6601_ (.A(net38),
    .B(_2220_),
    .COUT(_2221_),
    .SUM(_2222_));
 sky130_fd_sc_hd__ha_1 _6602_ (.A(net38),
    .B(net54),
    .COUT(_2223_),
    .SUM(_2224_));
 sky130_fd_sc_hd__ha_1 _6603_ (.A(_2090_),
    .B(net172),
    .COUT(_2225_),
    .SUM(_2226_));
 sky130_fd_sc_hd__ha_1 _6604_ (.A(_2227_),
    .B(_2228_),
    .COUT(_2229_),
    .SUM(_2230_));
 sky130_fd_sc_hd__ha_1 _6605_ (.A(_2105_),
    .B(_2231_),
    .COUT(_2232_),
    .SUM(_2233_));
 sky130_fd_sc_hd__ha_1 _6606_ (.A(_2234_),
    .B(_2207_),
    .COUT(_2235_),
    .SUM(_2236_));
 sky130_fd_sc_hd__ha_1 _6607_ (.A(_2237_),
    .B(_2208_),
    .COUT(_2116_),
    .SUM(_2238_));
 sky130_fd_sc_hd__ha_2 _6608_ (.A(_2239_),
    .B(net57),
    .COUT(_2240_),
    .SUM(_2241_));
 sky130_fd_sc_hd__ha_2 _6609_ (.A(net41),
    .B(_2242_),
    .COUT(_2243_),
    .SUM(_2244_));
 sky130_fd_sc_hd__ha_1 _6610_ (.A(net41),
    .B(net57),
    .COUT(_2245_),
    .SUM(_2246_));
 sky130_fd_sc_hd__ha_2 _6611_ (.A(_2247_),
    .B(net56),
    .COUT(_2248_),
    .SUM(_2249_));
 sky130_fd_sc_hd__ha_1 _6612_ (.A(net40),
    .B(_2250_),
    .COUT(_2251_),
    .SUM(_2252_));
 sky130_fd_sc_hd__ha_1 _6613_ (.A(net40),
    .B(net56),
    .COUT(_2253_),
    .SUM(_2254_));
 sky130_fd_sc_hd__ha_1 _6614_ (.A(_2255_),
    .B(net58),
    .COUT(_2256_),
    .SUM(_2257_));
 sky130_fd_sc_hd__ha_2 _6615_ (.A(net42),
    .B(_2258_),
    .COUT(_2259_),
    .SUM(_2260_));
 sky130_fd_sc_hd__ha_2 _6616_ (.A(net42),
    .B(net58),
    .COUT(_2261_),
    .SUM(_2262_));
 sky130_fd_sc_hd__ha_1 _6617_ (.A(_2263_),
    .B(_2264_),
    .COUT(_2265_),
    .SUM(_2266_));
 sky130_fd_sc_hd__ha_1 _6618_ (.A(_2267_),
    .B(_2268_),
    .COUT(_2269_),
    .SUM(_2270_));
 sky130_fd_sc_hd__ha_1 _6619_ (.A(_2271_),
    .B(_2272_),
    .COUT(_2273_),
    .SUM(_2274_));
 sky130_fd_sc_hd__ha_1 _6620_ (.A(_2275_),
    .B(_2276_),
    .COUT(_2277_),
    .SUM(_2278_));
 sky130_fd_sc_hd__ha_1 _6621_ (.A(_2279_),
    .B(_2096_),
    .COUT(_2280_),
    .SUM(_2281_));
 sky130_fd_sc_hd__ha_1 _6622_ (.A(_2100_),
    .B(_2101_),
    .COUT(_2282_),
    .SUM(_2283_));
 sky130_fd_sc_hd__ha_1 _6623_ (.A(net5),
    .B(_2284_),
    .COUT(_2285_),
    .SUM(_2286_));
 sky130_fd_sc_hd__ha_1 _6624_ (.A(_2287_),
    .B(_2111_),
    .COUT(_2288_),
    .SUM(_2289_));
 sky130_fd_sc_hd__ha_1 _6625_ (.A(_2290_),
    .B(net5),
    .COUT(_2291_),
    .SUM(_2292_));
 sky130_fd_sc_hd__ha_1 _6626_ (.A(_2293_),
    .B(_2092_),
    .COUT(_2294_),
    .SUM(_2295_));
 sky130_fd_sc_hd__ha_1 _6627_ (.A(_2296_),
    .B(_2111_),
    .COUT(_2297_),
    .SUM(_2298_));
 sky130_fd_sc_hd__ha_1 _6628_ (.A(_2299_),
    .B(_2092_),
    .COUT(_2300_),
    .SUM(_2301_));
 sky130_fd_sc_hd__ha_4 _6629_ (.A(_2111_),
    .B(_2302_),
    .COUT(_2303_),
    .SUM(_2304_));
 sky130_fd_sc_hd__ha_1 _6630_ (.A(_2305_),
    .B(_2111_),
    .COUT(_2306_),
    .SUM(_2307_));
 sky130_fd_sc_hd__ha_1 _6631_ (.A(_2308_),
    .B(_2111_),
    .COUT(_2309_),
    .SUM(_2310_));
 sky130_fd_sc_hd__ha_4 _6632_ (.A(_2311_),
    .B(_2092_),
    .COUT(_2312_),
    .SUM(_2313_));
 sky130_fd_sc_hd__ha_1 _6633_ (.A(_2107_),
    .B(_2092_),
    .COUT(_2314_),
    .SUM(_2315_));
 sky130_fd_sc_hd__ha_2 _6634_ (.A(_2316_),
    .B(_2317_),
    .COUT(_2318_),
    .SUM(_2319_));
 sky130_fd_sc_hd__ha_1 _6635_ (.A(_2320_),
    .B(_2321_),
    .COUT(_2322_),
    .SUM(_2323_));
 sky130_fd_sc_hd__ha_1 _6636_ (.A(_2324_),
    .B(_2237_),
    .COUT(_2325_),
    .SUM(_2326_));
 sky130_fd_sc_hd__ha_1 _6637_ (.A(_2327_),
    .B(_2328_),
    .COUT(_2329_),
    .SUM(_2330_));
 sky130_fd_sc_hd__ha_1 _6638_ (.A(_2098_),
    .B(_2113_),
    .COUT(_2332_),
    .SUM(_2333_));
 sky130_fd_sc_hd__ha_1 _6639_ (.A(_2101_),
    .B(_2334_),
    .COUT(_2331_),
    .SUM(_2335_));
 sky130_fd_sc_hd__ha_1 _6640_ (.A(_2336_),
    .B(_2238_),
    .COUT(_2337_),
    .SUM(_2338_));
 sky130_fd_sc_hd__ha_1 _6641_ (.A(_2339_),
    .B(net59),
    .COUT(_2340_),
    .SUM(_2341_));
 sky130_fd_sc_hd__ha_1 _6642_ (.A(net43),
    .B(_2342_),
    .COUT(_2343_),
    .SUM(_2344_));
 sky130_fd_sc_hd__ha_2 _6643_ (.A(net43),
    .B(net59),
    .COUT(_2345_),
    .SUM(_2346_));
 sky130_fd_sc_hd__ha_1 _6644_ (.A(_2347_),
    .B(net60),
    .COUT(_2348_),
    .SUM(_2349_));
 sky130_fd_sc_hd__ha_1 _6645_ (.A(net44),
    .B(_2350_),
    .COUT(_2351_),
    .SUM(_2352_));
 sky130_fd_sc_hd__ha_1 _6646_ (.A(net44),
    .B(net60),
    .COUT(_2353_),
    .SUM(_2354_));
 sky130_fd_sc_hd__ha_1 _6647_ (.A(_2355_),
    .B(_2356_),
    .COUT(_2357_),
    .SUM(_2358_));
 sky130_fd_sc_hd__ha_1 _6648_ (.A(_2359_),
    .B(_2360_),
    .COUT(_2361_),
    .SUM(_2362_));
 sky130_fd_sc_hd__ha_1 _6649_ (.A(_2363_),
    .B(net47),
    .COUT(_2364_),
    .SUM(_2365_));
 sky130_fd_sc_hd__ha_1 _6650_ (.A(net31),
    .B(_2366_),
    .COUT(_2367_),
    .SUM(_2368_));
 sky130_fd_sc_hd__ha_2 _6651_ (.A(net31),
    .B(net47),
    .COUT(_2369_),
    .SUM(_2370_));
 sky130_fd_sc_hd__ha_2 _6652_ (.A(_2371_),
    .B(net61),
    .COUT(_2372_),
    .SUM(_2373_));
 sky130_fd_sc_hd__ha_1 _6653_ (.A(net45),
    .B(_2374_),
    .COUT(_2375_),
    .SUM(_2376_));
 sky130_fd_sc_hd__ha_1 _6654_ (.A(net45),
    .B(net61),
    .COUT(_2377_),
    .SUM(_2378_));
 sky130_fd_sc_hd__ha_1 _6655_ (.A(_2379_),
    .B(_2380_),
    .COUT(_2381_),
    .SUM(_2382_));
 sky130_fd_sc_hd__ha_2 _6656_ (.A(_2383_),
    .B(_2384_),
    .COUT(_2385_),
    .SUM(_2386_));
 sky130_fd_sc_hd__ha_2 _6657_ (.A(_2387_),
    .B(_2388_),
    .COUT(_2389_),
    .SUM(_2390_));
 sky130_fd_sc_hd__ha_2 _6658_ (.A(_2391_),
    .B(_2392_),
    .COUT(_2393_),
    .SUM(_2394_));
 sky130_fd_sc_hd__ha_2 _6659_ (.A(_2395_),
    .B(_2396_),
    .COUT(_2397_),
    .SUM(_2398_));
 sky130_fd_sc_hd__ha_1 _6660_ (.A(_2399_),
    .B(_2400_),
    .COUT(_2401_),
    .SUM(_2402_));
 sky130_fd_sc_hd__ha_1 _6661_ (.A(_2403_),
    .B(_2404_),
    .COUT(_2405_),
    .SUM(_2406_));
 sky130_fd_sc_hd__ha_1 _6662_ (.A(_2407_),
    .B(_2408_),
    .COUT(_2409_),
    .SUM(_2410_));
 sky130_fd_sc_hd__ha_1 _6663_ (.A(_2411_),
    .B(_2412_),
    .COUT(_2413_),
    .SUM(_2414_));
 sky130_fd_sc_hd__ha_1 _6664_ (.A(_2415_),
    .B(_2416_),
    .COUT(_2417_),
    .SUM(_2418_));
 sky130_fd_sc_hd__ha_1 _6665_ (.A(_2419_),
    .B(_2420_),
    .COUT(_2421_),
    .SUM(_2422_));
 sky130_fd_sc_hd__ha_1 _6666_ (.A(_2423_),
    .B(_2424_),
    .COUT(_2425_),
    .SUM(_2426_));
 sky130_fd_sc_hd__ha_1 _6667_ (.A(_2427_),
    .B(_2428_),
    .COUT(_2429_),
    .SUM(_2430_));
 sky130_fd_sc_hd__ha_1 _6668_ (.A(_2121_),
    .B(_2103_),
    .COUT(_2431_),
    .SUM(_2432_));
 sky130_fd_sc_hd__ha_1 _6669_ (.A(_2433_),
    .B(_2124_),
    .COUT(_2434_),
    .SUM(_2435_));
 sky130_fd_sc_hd__ha_1 _6670_ (.A(_2436_),
    .B(_2124_),
    .COUT(_2437_),
    .SUM(_2438_));
 sky130_fd_sc_hd__ha_2 _6671_ (.A(_2439_),
    .B(_2124_),
    .COUT(_2440_),
    .SUM(_2441_));
 sky130_fd_sc_hd__ha_1 _6672_ (.A(_2442_),
    .B(net15),
    .COUT(_2444_),
    .SUM(_2445_));
 sky130_fd_sc_hd__ha_1 _6673_ (.A(_2446_),
    .B(_2124_),
    .COUT(_2447_),
    .SUM(_2448_));
 sky130_fd_sc_hd__ha_1 _6674_ (.A(_2449_),
    .B(_2124_),
    .COUT(_2450_),
    .SUM(_2451_));
 sky130_fd_sc_hd__ha_1 _6675_ (.A(_2452_),
    .B(net15),
    .COUT(_2453_),
    .SUM(_2454_));
 sky130_fd_sc_hd__ha_1 _6676_ (.A(_2455_),
    .B(net15),
    .COUT(_2456_),
    .SUM(_2457_));
 sky130_fd_sc_hd__ha_1 _6677_ (.A(_2458_),
    .B(_2443_),
    .COUT(_2459_),
    .SUM(_2460_));
 sky130_fd_sc_hd__ha_1 _6678_ (.A(_2461_),
    .B(_2443_),
    .COUT(_2462_),
    .SUM(_2463_));
 sky130_fd_sc_hd__ha_1 _6679_ (.A(_2464_),
    .B(_2443_),
    .COUT(_2465_),
    .SUM(_2466_));
 sky130_fd_sc_hd__ha_1 _6680_ (.A(_2109_),
    .B(_2443_),
    .COUT(_2467_),
    .SUM(_2468_));
 sky130_fd_sc_hd__ha_4 _6681_ (.A(_2124_),
    .B(_2110_),
    .COUT(_2469_),
    .SUM(_2470_));
 sky130_fd_sc_hd__ha_4 _6682_ (.A(_2471_),
    .B(_2122_),
    .COUT(_2472_),
    .SUM(_2473_));
 sky130_fd_sc_hd__ha_4 _6683_ (.A(_2474_),
    .B(_2443_),
    .COUT(_2475_),
    .SUM(_2476_));
 sky130_fd_sc_hd__ha_1 _6684_ (.A(_2477_),
    .B(_2478_),
    .COUT(_2479_),
    .SUM(_2480_));
 sky130_fd_sc_hd__ha_1 _6685_ (.A(_2481_),
    .B(_2482_),
    .COUT(_2483_),
    .SUM(_2484_));
 sky130_fd_sc_hd__ha_1 _6686_ (.A(_2485_),
    .B(_2336_),
    .COUT(_2486_),
    .SUM(_2487_));
 sky130_fd_sc_hd__ha_1 _6687_ (.A(_2488_),
    .B(_2489_),
    .COUT(_2490_),
    .SUM(_2491_));
 sky130_fd_sc_hd__ha_1 _6688_ (.A(_2492_),
    .B(_2493_),
    .COUT(_2494_),
    .SUM(_2495_));
 sky130_fd_sc_hd__ha_1 _6689_ (.A(_2115_),
    .B(_2128_),
    .COUT(_2496_),
    .SUM(_2497_));
 sky130_fd_sc_hd__ha_1 _6690_ (.A(_2335_),
    .B(_2424_),
    .COUT(_2112_),
    .SUM(_2498_));
 sky130_fd_sc_hd__ha_1 _6691_ (.A(_2499_),
    .B(_2338_),
    .COUT(_2140_),
    .SUM(_2500_));
 sky130_fd_sc_hd__ha_1 _6692_ (.A(_2501_),
    .B(_2502_),
    .COUT(_2503_),
    .SUM(_2504_));
 sky130_fd_sc_hd__ha_2 _6693_ (.A(_2505_),
    .B(_2506_),
    .COUT(_2507_),
    .SUM(_2508_));
 sky130_fd_sc_hd__ha_1 _6694_ (.A(_2509_),
    .B(net49),
    .COUT(_2510_),
    .SUM(_2511_));
 sky130_fd_sc_hd__ha_1 _6695_ (.A(net33),
    .B(_2512_),
    .COUT(_2513_),
    .SUM(_2514_));
 sky130_fd_sc_hd__ha_1 _6696_ (.A(net33),
    .B(net49),
    .COUT(_2515_),
    .SUM(_2516_));
 sky130_fd_sc_hd__ha_1 _6697_ (.A(_2517_),
    .B(net48),
    .COUT(_2518_),
    .SUM(_2519_));
 sky130_fd_sc_hd__ha_1 _6698_ (.A(net32),
    .B(_2520_),
    .COUT(_2521_),
    .SUM(_2522_));
 sky130_fd_sc_hd__ha_1 _6699_ (.A(net32),
    .B(net48),
    .COUT(_2523_),
    .SUM(_2524_));
 sky130_fd_sc_hd__ha_1 _6700_ (.A(_2525_),
    .B(_2526_),
    .COUT(_2527_),
    .SUM(_2528_));
 sky130_fd_sc_hd__ha_1 _6701_ (.A(_2529_),
    .B(_2530_),
    .COUT(_2531_),
    .SUM(_2532_));
 sky130_fd_sc_hd__ha_1 _6702_ (.A(_2533_),
    .B(_2534_),
    .COUT(_2535_),
    .SUM(_2536_));
 sky130_fd_sc_hd__ha_1 _6703_ (.A(_2537_),
    .B(_2538_),
    .COUT(_2539_),
    .SUM(_2540_));
 sky130_fd_sc_hd__ha_1 _6704_ (.A(_2541_),
    .B(net51),
    .COUT(_2542_),
    .SUM(_2543_));
 sky130_fd_sc_hd__ha_1 _6705_ (.A(net35),
    .B(_2544_),
    .COUT(_2545_),
    .SUM(_2546_));
 sky130_fd_sc_hd__ha_1 _6706_ (.A(net35),
    .B(net51),
    .COUT(_2547_),
    .SUM(_2548_));
 sky130_fd_sc_hd__ha_2 _6707_ (.A(_2549_),
    .B(net50),
    .COUT(_2550_),
    .SUM(_2551_));
 sky130_fd_sc_hd__ha_1 _6708_ (.A(net34),
    .B(_2552_),
    .COUT(_2553_),
    .SUM(_2554_));
 sky130_fd_sc_hd__ha_1 _6709_ (.A(net34),
    .B(net50),
    .COUT(_2555_),
    .SUM(_2556_));
 sky130_fd_sc_hd__ha_1 _6710_ (.A(_2557_),
    .B(_2558_),
    .COUT(_2559_),
    .SUM(_2560_));
 sky130_fd_sc_hd__ha_1 _6711_ (.A(_2561_),
    .B(_2562_),
    .COUT(_2563_),
    .SUM(_2564_));
 sky130_fd_sc_hd__ha_1 _6712_ (.A(_2565_),
    .B(_2566_),
    .COUT(_2567_),
    .SUM(_2568_));
 sky130_fd_sc_hd__ha_1 _6713_ (.A(_2569_),
    .B(_2570_),
    .COUT(_2571_),
    .SUM(_2572_));
 sky130_fd_sc_hd__ha_2 _6714_ (.A(_2573_),
    .B(_2574_),
    .COUT(_2575_),
    .SUM(_2576_));
 sky130_fd_sc_hd__ha_1 _6715_ (.A(_2577_),
    .B(_2578_),
    .COUT(_2579_),
    .SUM(_2580_));
 sky130_fd_sc_hd__ha_1 _6716_ (.A(_2581_),
    .B(_2582_),
    .COUT(_2583_),
    .SUM(_2584_));
 sky130_fd_sc_hd__ha_1 _6717_ (.A(_2585_),
    .B(_2586_),
    .COUT(_2587_),
    .SUM(_2588_));
 sky130_fd_sc_hd__ha_2 _6718_ (.A(_2589_),
    .B(_2590_),
    .COUT(_2591_),
    .SUM(_2592_));
 sky130_fd_sc_hd__ha_2 _6719_ (.A(_2593_),
    .B(_2594_),
    .COUT(_2595_),
    .SUM(_2596_));
 sky130_fd_sc_hd__ha_2 _6720_ (.A(_2597_),
    .B(_2598_),
    .COUT(_2599_),
    .SUM(_2600_));
 sky130_fd_sc_hd__ha_2 _6721_ (.A(_2601_),
    .B(_2602_),
    .COUT(_2603_),
    .SUM(_2604_));
 sky130_fd_sc_hd__ha_2 _6722_ (.A(_2605_),
    .B(_2606_),
    .COUT(_2607_),
    .SUM(_2608_));
 sky130_fd_sc_hd__ha_1 _6723_ (.A(_2609_),
    .B(_2610_),
    .COUT(_2611_),
    .SUM(_2612_));
 sky130_fd_sc_hd__ha_1 _6724_ (.A(_2613_),
    .B(_2614_),
    .COUT(_2615_),
    .SUM(_2616_));
 sky130_fd_sc_hd__ha_1 _6725_ (.A(_2617_),
    .B(_2618_),
    .COUT(_2619_),
    .SUM(_2620_));
 sky130_fd_sc_hd__ha_2 _6726_ (.A(_2621_),
    .B(_2622_),
    .COUT(_2623_),
    .SUM(_2624_));
 sky130_fd_sc_hd__ha_1 _6727_ (.A(_2625_),
    .B(_2626_),
    .COUT(_2627_),
    .SUM(_2628_));
 sky130_fd_sc_hd__ha_1 _6728_ (.A(_2629_),
    .B(_2630_),
    .COUT(_2631_),
    .SUM(_2632_));
 sky130_fd_sc_hd__ha_1 _6729_ (.A(_2633_),
    .B(_2634_),
    .COUT(_2635_),
    .SUM(_2636_));
 sky130_fd_sc_hd__ha_1 _6730_ (.A(_2637_),
    .B(_2638_),
    .COUT(_2639_),
    .SUM(_2640_));
 sky130_fd_sc_hd__ha_1 _6731_ (.A(_2641_),
    .B(_2642_),
    .COUT(_2643_),
    .SUM(_2644_));
 sky130_fd_sc_hd__ha_1 _6732_ (.A(_2645_),
    .B(_2646_),
    .COUT(_2647_),
    .SUM(_2648_));
 sky130_fd_sc_hd__ha_1 _6733_ (.A(_2132_),
    .B(_2133_),
    .COUT(_2649_),
    .SUM(_2650_));
 sky130_fd_sc_hd__ha_1 _6734_ (.A(_2651_),
    .B(net14),
    .COUT(_2653_),
    .SUM(_2654_));
 sky130_fd_sc_hd__ha_1 _6735_ (.A(_2655_),
    .B(net14),
    .COUT(_2656_),
    .SUM(_2657_));
 sky130_fd_sc_hd__ha_1 _6736_ (.A(_2658_),
    .B(net9),
    .COUT(_2659_),
    .SUM(_2660_));
 sky130_fd_sc_hd__ha_1 _6737_ (.A(_2661_),
    .B(net14),
    .COUT(_2662_),
    .SUM(_2663_));
 sky130_fd_sc_hd__ha_1 _6738_ (.A(_2664_),
    .B(_2665_),
    .COUT(_2666_),
    .SUM(_2667_));
 sky130_fd_sc_hd__ha_1 _6739_ (.A(_2668_),
    .B(net14),
    .COUT(_2669_),
    .SUM(_2670_));
 sky130_fd_sc_hd__ha_1 _6740_ (.A(_2671_),
    .B(_2665_),
    .COUT(_2672_),
    .SUM(_2673_));
 sky130_fd_sc_hd__ha_1 _6741_ (.A(_2674_),
    .B(net14),
    .COUT(_2675_),
    .SUM(_2676_));
 sky130_fd_sc_hd__ha_1 _6742_ (.A(_2677_),
    .B(_2652_),
    .COUT(_2678_),
    .SUM(_2679_));
 sky130_fd_sc_hd__ha_1 _6743_ (.A(_2680_),
    .B(_2652_),
    .COUT(_2681_),
    .SUM(_2682_));
 sky130_fd_sc_hd__ha_1 _6744_ (.A(_2683_),
    .B(_2665_),
    .COUT(_2684_),
    .SUM(_2685_));
 sky130_fd_sc_hd__ha_1 _6745_ (.A(_2686_),
    .B(_2652_),
    .COUT(_2687_),
    .SUM(_2688_));
 sky130_fd_sc_hd__ha_1 _6746_ (.A(_2689_),
    .B(_2652_),
    .COUT(_2690_),
    .SUM(_2691_));
 sky130_fd_sc_hd__ha_4 _6747_ (.A(_2692_),
    .B(_2652_),
    .COUT(_2693_),
    .SUM(_2694_));
 sky130_fd_sc_hd__ha_1 _6748_ (.A(_2695_),
    .B(_2696_),
    .COUT(_2697_),
    .SUM(_2698_));
 sky130_fd_sc_hd__ha_1 _6749_ (.A(_2699_),
    .B(_2700_),
    .COUT(_2701_),
    .SUM(_2702_));
 sky130_fd_sc_hd__ha_1 _6750_ (.A(_2703_),
    .B(_2499_),
    .COUT(_2704_),
    .SUM(_2705_));
 sky130_fd_sc_hd__ha_1 _6751_ (.A(_2706_),
    .B(_2707_),
    .COUT(_2708_),
    .SUM(_2709_));
 sky130_fd_sc_hd__ha_1 _6752_ (.A(_2710_),
    .B(_2711_),
    .COUT(_2712_),
    .SUM(_2713_));
 sky130_fd_sc_hd__ha_1 _6753_ (.A(_2714_),
    .B(_2715_),
    .COUT(_2716_),
    .SUM(_2717_));
 sky130_fd_sc_hd__ha_1 _6754_ (.A(_2130_),
    .B(_2137_),
    .COUT(_2718_),
    .SUM(_2719_));
 sky130_fd_sc_hd__ha_1 _6755_ (.A(_2498_),
    .B(_2638_),
    .COUT(_2127_),
    .SUM(_2720_));
 sky130_fd_sc_hd__ha_1 _6756_ (.A(_2721_),
    .B(_2500_),
    .COUT(_2150_),
    .SUM(_2722_));
 sky130_fd_sc_hd__ha_1 _6757_ (.A(_2723_),
    .B(_2724_),
    .COUT(_2725_),
    .SUM(_2726_));
 sky130_fd_sc_hd__ha_2 _6758_ (.A(_2727_),
    .B(_2728_),
    .COUT(_2729_),
    .SUM(_2730_));
 sky130_fd_sc_hd__ha_1 _6759_ (.A(_2731_),
    .B(_2732_),
    .COUT(_2733_),
    .SUM(_2734_));
 sky130_fd_sc_hd__ha_2 _6760_ (.A(_2735_),
    .B(_2736_),
    .COUT(_2737_),
    .SUM(_2738_));
 sky130_fd_sc_hd__ha_2 _6761_ (.A(_2739_),
    .B(_2740_),
    .COUT(_2741_),
    .SUM(_2742_));
 sky130_fd_sc_hd__ha_2 _6762_ (.A(_2743_),
    .B(_2744_),
    .COUT(_2745_),
    .SUM(_2746_));
 sky130_fd_sc_hd__ha_1 _6763_ (.A(_2747_),
    .B(_2748_),
    .COUT(_2749_),
    .SUM(_2750_));
 sky130_fd_sc_hd__ha_2 _6764_ (.A(_2751_),
    .B(_2752_),
    .COUT(_2753_),
    .SUM(_2754_));
 sky130_fd_sc_hd__ha_2 _6765_ (.A(_2755_),
    .B(_2756_),
    .COUT(_2757_),
    .SUM(_2758_));
 sky130_fd_sc_hd__ha_1 _6766_ (.A(_2759_),
    .B(_2760_),
    .COUT(_2761_),
    .SUM(_2762_));
 sky130_fd_sc_hd__ha_2 _6767_ (.A(_2763_),
    .B(_2764_),
    .COUT(_2765_),
    .SUM(_2766_));
 sky130_fd_sc_hd__ha_1 _6768_ (.A(_2767_),
    .B(_2768_),
    .COUT(_2769_),
    .SUM(_2770_));
 sky130_fd_sc_hd__ha_1 _6769_ (.A(_2771_),
    .B(_2772_),
    .COUT(_2773_),
    .SUM(_2774_));
 sky130_fd_sc_hd__ha_2 _6770_ (.A(_2771_),
    .B(_2772_),
    .COUT(_2775_),
    .SUM(_2776_));
 sky130_fd_sc_hd__ha_1 _6771_ (.A(_2777_),
    .B(_2778_),
    .COUT(_2779_),
    .SUM(_2780_));
 sky130_fd_sc_hd__ha_1 _6772_ (.A(_2781_),
    .B(_2782_),
    .COUT(_2783_),
    .SUM(_2784_));
 sky130_fd_sc_hd__ha_1 _6773_ (.A(_2785_),
    .B(_2786_),
    .COUT(_2787_),
    .SUM(_2788_));
 sky130_fd_sc_hd__ha_1 _6774_ (.A(_2789_),
    .B(_2790_),
    .COUT(_2791_),
    .SUM(_2792_));
 sky130_fd_sc_hd__ha_1 _6775_ (.A(_2793_),
    .B(_2794_),
    .COUT(_2795_),
    .SUM(_2796_));
 sky130_fd_sc_hd__ha_1 _6776_ (.A(_2797_),
    .B(_2798_),
    .COUT(_2799_),
    .SUM(_2800_));
 sky130_fd_sc_hd__ha_1 _6777_ (.A(_2801_),
    .B(_2802_),
    .COUT(_2803_),
    .SUM(_2804_));
 sky130_fd_sc_hd__ha_2 _6778_ (.A(_2805_),
    .B(_2806_),
    .COUT(_2807_),
    .SUM(_2808_));
 sky130_fd_sc_hd__ha_1 _6779_ (.A(_2809_),
    .B(_2810_),
    .COUT(_2811_),
    .SUM(_2812_));
 sky130_fd_sc_hd__ha_1 _6780_ (.A(_2813_),
    .B(_2814_),
    .COUT(_2815_),
    .SUM(_2816_));
 sky130_fd_sc_hd__ha_1 _6781_ (.A(_2817_),
    .B(_2818_),
    .COUT(_2819_),
    .SUM(_2820_));
 sky130_fd_sc_hd__ha_1 _6782_ (.A(_2821_),
    .B(_2822_),
    .COUT(_2823_),
    .SUM(_2824_));
 sky130_fd_sc_hd__ha_1 _6783_ (.A(_2825_),
    .B(_2826_),
    .COUT(_2827_),
    .SUM(_2828_));
 sky130_fd_sc_hd__ha_1 _6784_ (.A(_2829_),
    .B(_2830_),
    .COUT(_2831_),
    .SUM(_2832_));
 sky130_fd_sc_hd__ha_1 _6785_ (.A(_2833_),
    .B(_2834_),
    .COUT(_2835_),
    .SUM(_2836_));
 sky130_fd_sc_hd__ha_1 _6786_ (.A(_2837_),
    .B(_2838_),
    .COUT(_2839_),
    .SUM(_2840_));
 sky130_fd_sc_hd__ha_1 _6787_ (.A(_2841_),
    .B(_2842_),
    .COUT(_2843_),
    .SUM(_2844_));
 sky130_fd_sc_hd__ha_1 _6788_ (.A(_2145_),
    .B(_2135_),
    .COUT(_2845_),
    .SUM(_2846_));
 sky130_fd_sc_hd__ha_1 _6789_ (.A(_2847_),
    .B(_2848_),
    .COUT(_2849_),
    .SUM(_2850_));
 sky130_fd_sc_hd__ha_1 _6790_ (.A(_2851_),
    .B(net12),
    .COUT(_2853_),
    .SUM(_2854_));
 sky130_fd_sc_hd__ha_1 _6791_ (.A(_2855_),
    .B(net12),
    .COUT(_2856_),
    .SUM(_2857_));
 sky130_fd_sc_hd__ha_1 _6792_ (.A(_2858_),
    .B(_2852_),
    .COUT(_2859_),
    .SUM(_2860_));
 sky130_fd_sc_hd__ha_1 _6793_ (.A(_2861_),
    .B(_2852_),
    .COUT(_2862_),
    .SUM(_2863_));
 sky130_fd_sc_hd__ha_1 _6794_ (.A(_2864_),
    .B(_2852_),
    .COUT(_2865_),
    .SUM(_2866_));
 sky130_fd_sc_hd__ha_1 _6795_ (.A(_2867_),
    .B(_2868_),
    .COUT(_2869_),
    .SUM(_2870_));
 sky130_fd_sc_hd__ha_1 _6796_ (.A(_2871_),
    .B(_2852_),
    .COUT(_2872_),
    .SUM(_2873_));
 sky130_fd_sc_hd__ha_1 _6797_ (.A(_2874_),
    .B(_2868_),
    .COUT(_2875_),
    .SUM(_2876_));
 sky130_fd_sc_hd__ha_1 _6798_ (.A(_2877_),
    .B(_2852_),
    .COUT(_2878_),
    .SUM(_2879_));
 sky130_fd_sc_hd__ha_1 _6799_ (.A(_2880_),
    .B(_2852_),
    .COUT(_2881_),
    .SUM(_2882_));
 sky130_fd_sc_hd__ha_1 _6800_ (.A(_2883_),
    .B(_2852_),
    .COUT(_2884_),
    .SUM(_2885_));
 sky130_fd_sc_hd__ha_1 _6801_ (.A(_2886_),
    .B(_2868_),
    .COUT(_2887_),
    .SUM(_2888_));
 sky130_fd_sc_hd__ha_4 _6802_ (.A(_2889_),
    .B(_2852_),
    .COUT(_2890_),
    .SUM(_2891_));
 sky130_fd_sc_hd__ha_4 _6803_ (.A(_2892_),
    .B(_2868_),
    .COUT(_2893_),
    .SUM(_2894_));
 sky130_fd_sc_hd__ha_1 _6804_ (.A(_2895_),
    .B(_2896_),
    .COUT(_2897_),
    .SUM(_2898_));
 sky130_fd_sc_hd__ha_2 _6805_ (.A(_2899_),
    .B(_2900_),
    .COUT(_2901_),
    .SUM(_2902_));
 sky130_fd_sc_hd__ha_1 _6806_ (.A(_2903_),
    .B(_2721_),
    .COUT(_2904_),
    .SUM(_2905_));
 sky130_fd_sc_hd__ha_1 _6807_ (.A(_2906_),
    .B(_2907_),
    .COUT(_2908_),
    .SUM(_2909_));
 sky130_fd_sc_hd__ha_1 _6808_ (.A(_2910_),
    .B(_2911_),
    .COUT(_2912_),
    .SUM(_2913_));
 sky130_fd_sc_hd__ha_1 _6809_ (.A(_2914_),
    .B(_2915_),
    .COUT(_2916_),
    .SUM(_2917_));
 sky130_fd_sc_hd__ha_1 _6810_ (.A(_2918_),
    .B(_2919_),
    .COUT(_2920_),
    .SUM(_2921_));
 sky130_fd_sc_hd__ha_1 _6811_ (.A(_2139_),
    .B(_2147_),
    .COUT(_2922_),
    .SUM(_2923_));
 sky130_fd_sc_hd__ha_1 _6812_ (.A(_2720_),
    .B(_2830_),
    .COUT(_2136_),
    .SUM(_2924_));
 sky130_fd_sc_hd__ha_1 _6813_ (.A(_2925_),
    .B(_2722_),
    .COUT(_2165_),
    .SUM(_2926_));
 sky130_fd_sc_hd__ha_1 _6814_ (.A(_2927_),
    .B(_2928_),
    .COUT(_2929_),
    .SUM(_2930_));
 sky130_fd_sc_hd__ha_1 _6815_ (.A(_2931_),
    .B(_2932_),
    .COUT(_2933_),
    .SUM(_2934_));
 sky130_fd_sc_hd__ha_2 _6816_ (.A(_2935_),
    .B(_2936_),
    .COUT(_2937_),
    .SUM(_2938_));
 sky130_fd_sc_hd__ha_2 _6817_ (.A(_2939_),
    .B(_2940_),
    .COUT(_2941_),
    .SUM(_2942_));
 sky130_fd_sc_hd__ha_1 _6818_ (.A(_2943_),
    .B(_2944_),
    .COUT(_2945_),
    .SUM(_2946_));
 sky130_fd_sc_hd__ha_2 _6819_ (.A(_2947_),
    .B(_2948_),
    .COUT(_2949_),
    .SUM(_2950_));
 sky130_fd_sc_hd__ha_1 _6820_ (.A(_2951_),
    .B(_2952_),
    .COUT(_2953_),
    .SUM(_2954_));
 sky130_fd_sc_hd__ha_2 _6821_ (.A(_2951_),
    .B(_2952_),
    .COUT(_2955_),
    .SUM(_2956_));
 sky130_fd_sc_hd__ha_2 _6822_ (.A(_2957_),
    .B(_2958_),
    .COUT(_2959_),
    .SUM(_2960_));
 sky130_fd_sc_hd__ha_1 _6823_ (.A(_2961_),
    .B(_2962_),
    .COUT(_2963_),
    .SUM(_2964_));
 sky130_fd_sc_hd__ha_1 _6824_ (.A(_2965_),
    .B(_2966_),
    .COUT(_2967_),
    .SUM(_2968_));
 sky130_fd_sc_hd__ha_2 _6825_ (.A(_2969_),
    .B(_2970_),
    .COUT(_2971_),
    .SUM(_2972_));
 sky130_fd_sc_hd__ha_2 _6826_ (.A(_2973_),
    .B(_2974_),
    .COUT(_2975_),
    .SUM(_2976_));
 sky130_fd_sc_hd__ha_2 _6827_ (.A(_2977_),
    .B(_2978_),
    .COUT(_2979_),
    .SUM(_2980_));
 sky130_fd_sc_hd__ha_1 _6828_ (.A(_2981_),
    .B(_2982_),
    .COUT(_2983_),
    .SUM(_2984_));
 sky130_fd_sc_hd__ha_1 _6829_ (.A(_2985_),
    .B(_2986_),
    .COUT(_2987_),
    .SUM(_2988_));
 sky130_fd_sc_hd__ha_1 _6830_ (.A(_2985_),
    .B(_2986_),
    .COUT(_2989_),
    .SUM(_2990_));
 sky130_fd_sc_hd__ha_1 _6831_ (.A(_2991_),
    .B(_2992_),
    .COUT(_2993_),
    .SUM(_2994_));
 sky130_fd_sc_hd__ha_2 _6832_ (.A(_2995_),
    .B(_2996_),
    .COUT(_2997_),
    .SUM(_2998_));
 sky130_fd_sc_hd__ha_1 _6833_ (.A(_2999_),
    .B(_3000_),
    .COUT(_3001_),
    .SUM(_3002_));
 sky130_fd_sc_hd__ha_2 _6834_ (.A(_3003_),
    .B(_3004_),
    .COUT(_3005_),
    .SUM(_3006_));
 sky130_fd_sc_hd__ha_1 _6835_ (.A(_3007_),
    .B(_3008_),
    .COUT(_3009_),
    .SUM(_3010_));
 sky130_fd_sc_hd__ha_1 _6836_ (.A(_3011_),
    .B(_3012_),
    .COUT(_3013_),
    .SUM(_3014_));
 sky130_fd_sc_hd__ha_1 _6837_ (.A(_3015_),
    .B(_3016_),
    .COUT(_3017_),
    .SUM(_3018_));
 sky130_fd_sc_hd__ha_1 _6838_ (.A(_3019_),
    .B(_3020_),
    .COUT(_3021_),
    .SUM(_3022_));
 sky130_fd_sc_hd__ha_1 _6839_ (.A(_3023_),
    .B(_3024_),
    .COUT(_3025_),
    .SUM(_3026_));
 sky130_fd_sc_hd__ha_1 _6840_ (.A(_2154_),
    .B(_2155_),
    .COUT(_3027_),
    .SUM(_3028_));
 sky130_fd_sc_hd__ha_1 _6841_ (.A(_3029_),
    .B(_3030_),
    .COUT(_3031_),
    .SUM(_3032_));
 sky130_fd_sc_hd__ha_2 _6842_ (.A(_3033_),
    .B(_3034_),
    .COUT(_3035_),
    .SUM(_3036_));
 sky130_fd_sc_hd__ha_1 _6843_ (.A(_3037_),
    .B(net24),
    .COUT(_3039_),
    .SUM(_3040_));
 sky130_fd_sc_hd__ha_1 _6844_ (.A(_3041_),
    .B(net24),
    .COUT(_3042_),
    .SUM(_3043_));
 sky130_fd_sc_hd__ha_1 _6845_ (.A(_3044_),
    .B(net24),
    .COUT(_3045_),
    .SUM(_3046_));
 sky130_fd_sc_hd__ha_1 _6846_ (.A(_3047_),
    .B(net24),
    .COUT(_3048_),
    .SUM(_3049_));
 sky130_fd_sc_hd__ha_1 _6847_ (.A(_3050_),
    .B(net24),
    .COUT(_3051_),
    .SUM(_3052_));
 sky130_fd_sc_hd__ha_1 _6848_ (.A(_3053_),
    .B(net26),
    .COUT(_3054_),
    .SUM(_3055_));
 sky130_fd_sc_hd__ha_1 _6849_ (.A(_3056_),
    .B(_3057_),
    .COUT(_3058_),
    .SUM(_3059_));
 sky130_fd_sc_hd__ha_1 _6850_ (.A(_3060_),
    .B(net26),
    .COUT(_3061_),
    .SUM(_3062_));
 sky130_fd_sc_hd__ha_1 _6851_ (.A(_3063_),
    .B(_3057_),
    .COUT(_3064_),
    .SUM(_3065_));
 sky130_fd_sc_hd__ha_1 _6852_ (.A(_3066_),
    .B(_3038_),
    .COUT(_3067_),
    .SUM(_3068_));
 sky130_fd_sc_hd__ha_1 _6853_ (.A(_3069_),
    .B(_3038_),
    .COUT(_3070_),
    .SUM(_3071_));
 sky130_fd_sc_hd__ha_1 _6854_ (.A(_3072_),
    .B(_3038_),
    .COUT(_3073_),
    .SUM(_3074_));
 sky130_fd_sc_hd__ha_1 _6855_ (.A(_3075_),
    .B(_3057_),
    .COUT(_3076_),
    .SUM(_3077_));
 sky130_fd_sc_hd__ha_4 _6856_ (.A(_3038_),
    .B(_3078_),
    .COUT(_3079_),
    .SUM(_3080_));
 sky130_fd_sc_hd__ha_1 _6857_ (.A(_3081_),
    .B(_3082_),
    .COUT(_3083_),
    .SUM(_3084_));
 sky130_fd_sc_hd__ha_1 _6858_ (.A(_3085_),
    .B(_3086_),
    .COUT(_3087_),
    .SUM(_3088_));
 sky130_fd_sc_hd__ha_1 _6859_ (.A(_3089_),
    .B(_2925_),
    .COUT(_3090_),
    .SUM(_3091_));
 sky130_fd_sc_hd__ha_1 _6860_ (.A(_3092_),
    .B(_3093_),
    .COUT(_3094_),
    .SUM(_3095_));
 sky130_fd_sc_hd__ha_1 _6861_ (.A(_3096_),
    .B(_3097_),
    .COUT(_3098_),
    .SUM(_3099_));
 sky130_fd_sc_hd__ha_1 _6862_ (.A(_3100_),
    .B(_3101_),
    .COUT(_3102_),
    .SUM(_3103_));
 sky130_fd_sc_hd__ha_1 _6863_ (.A(_3104_),
    .B(_3105_),
    .COUT(_3106_),
    .SUM(_3107_));
 sky130_fd_sc_hd__ha_1 _6864_ (.A(_3108_),
    .B(_3109_),
    .COUT(_3110_),
    .SUM(_3111_));
 sky130_fd_sc_hd__ha_1 _6865_ (.A(_2149_),
    .B(_2157_),
    .COUT(_3112_),
    .SUM(_3113_));
 sky130_fd_sc_hd__ha_1 _6866_ (.A(_2924_),
    .B(_3008_),
    .COUT(_2146_),
    .SUM(_3114_));
 sky130_fd_sc_hd__ha_1 _6867_ (.A(_3115_),
    .B(_2926_),
    .COUT(_2174_),
    .SUM(_3116_));
 sky130_fd_sc_hd__ha_2 _6868_ (.A(_3117_),
    .B(_3118_),
    .COUT(_3119_),
    .SUM(_3120_));
 sky130_fd_sc_hd__ha_1 _6869_ (.A(_3121_),
    .B(_3122_),
    .COUT(_3123_),
    .SUM(_3124_));
 sky130_fd_sc_hd__ha_2 _6870_ (.A(_3125_),
    .B(_3126_),
    .COUT(_3127_),
    .SUM(_3128_));
 sky130_fd_sc_hd__ha_1 _6871_ (.A(_3129_),
    .B(_3130_),
    .COUT(_3131_),
    .SUM(_3132_));
 sky130_fd_sc_hd__ha_1 _6872_ (.A(_3133_),
    .B(_3134_),
    .COUT(_3135_),
    .SUM(_3136_));
 sky130_fd_sc_hd__ha_1 _6873_ (.A(_3137_),
    .B(_3138_),
    .COUT(_3139_),
    .SUM(_3140_));
 sky130_fd_sc_hd__ha_1 _6874_ (.A(_3141_),
    .B(_3142_),
    .COUT(_3143_),
    .SUM(_3144_));
 sky130_fd_sc_hd__ha_1 _6875_ (.A(_3145_),
    .B(_3146_),
    .COUT(_3147_),
    .SUM(_3148_));
 sky130_fd_sc_hd__ha_2 _6876_ (.A(_3133_),
    .B(_3134_),
    .COUT(_3149_),
    .SUM(_3150_));
 sky130_fd_sc_hd__ha_1 _6877_ (.A(_3151_),
    .B(_3152_),
    .COUT(_3153_),
    .SUM(_3154_));
 sky130_fd_sc_hd__ha_1 _6878_ (.A(_3155_),
    .B(_3156_),
    .COUT(_3157_),
    .SUM(_3158_));
 sky130_fd_sc_hd__ha_1 _6879_ (.A(_3159_),
    .B(_3160_),
    .COUT(_3161_),
    .SUM(_3162_));
 sky130_fd_sc_hd__ha_1 _6880_ (.A(_3163_),
    .B(_3164_),
    .COUT(_3165_),
    .SUM(_3166_));
 sky130_fd_sc_hd__ha_1 _6881_ (.A(_3167_),
    .B(_3168_),
    .COUT(_3169_),
    .SUM(_3170_));
 sky130_fd_sc_hd__ha_1 _6882_ (.A(_3171_),
    .B(_3172_),
    .COUT(_3173_),
    .SUM(_3174_));
 sky130_fd_sc_hd__ha_1 _6883_ (.A(_3175_),
    .B(_3176_),
    .COUT(_3177_),
    .SUM(_3178_));
 sky130_fd_sc_hd__ha_1 _6884_ (.A(_3179_),
    .B(_3180_),
    .COUT(_3181_),
    .SUM(_3182_));
 sky130_fd_sc_hd__ha_1 _6885_ (.A(_3183_),
    .B(_3184_),
    .COUT(_3185_),
    .SUM(_3186_));
 sky130_fd_sc_hd__ha_1 _6886_ (.A(_3187_),
    .B(_3188_),
    .COUT(_3189_),
    .SUM(_3190_));
 sky130_fd_sc_hd__ha_1 _6887_ (.A(_3191_),
    .B(_3192_),
    .COUT(_3193_),
    .SUM(_3194_));
 sky130_fd_sc_hd__ha_1 _6888_ (.A(_2160_),
    .B(_2161_),
    .COUT(_3195_),
    .SUM(_3196_));
 sky130_fd_sc_hd__ha_2 _6889_ (.A(_3197_),
    .B(_3198_),
    .COUT(_3199_),
    .SUM(_3200_));
 sky130_fd_sc_hd__ha_1 _6890_ (.A(_3201_),
    .B(_3202_),
    .COUT(_3203_),
    .SUM(_3204_));
 sky130_fd_sc_hd__ha_2 _6891_ (.A(_3205_),
    .B(_3206_),
    .COUT(_3207_),
    .SUM(_3208_));
 sky130_fd_sc_hd__ha_2 _6892_ (.A(_3209_),
    .B(_3210_),
    .COUT(_3211_),
    .SUM(_3212_));
 sky130_fd_sc_hd__ha_1 _6893_ (.A(net10),
    .B(_3214_),
    .COUT(_3215_),
    .SUM(_3216_));
 sky130_fd_sc_hd__ha_1 _6894_ (.A(net10),
    .B(_3217_),
    .COUT(_3218_),
    .SUM(_3219_));
 sky130_fd_sc_hd__ha_1 _6895_ (.A(net10),
    .B(_3220_),
    .COUT(_3221_),
    .SUM(_3222_));
 sky130_fd_sc_hd__ha_1 _6896_ (.A(net10),
    .B(_3223_),
    .COUT(_3224_),
    .SUM(_3225_));
 sky130_fd_sc_hd__ha_1 _6897_ (.A(net10),
    .B(_3226_),
    .COUT(_3227_),
    .SUM(_3228_));
 sky130_fd_sc_hd__ha_1 _6898_ (.A(net10),
    .B(_3229_),
    .COUT(_3230_),
    .SUM(_3231_));
 sky130_fd_sc_hd__ha_1 _6899_ (.A(net19),
    .B(_3232_),
    .COUT(_3233_),
    .SUM(_3234_));
 sky130_fd_sc_hd__ha_1 _6900_ (.A(net11),
    .B(_3236_),
    .COUT(_3237_),
    .SUM(_3238_));
 sky130_fd_sc_hd__ha_1 _6901_ (.A(_3239_),
    .B(net19),
    .COUT(_3240_),
    .SUM(_3241_));
 sky130_fd_sc_hd__ha_1 _6902_ (.A(_3235_),
    .B(_3242_),
    .COUT(_3243_),
    .SUM(_3244_));
 sky130_fd_sc_hd__ha_1 _6903_ (.A(net19),
    .B(_3245_),
    .COUT(_3246_),
    .SUM(_3247_));
 sky130_fd_sc_hd__ha_1 _6904_ (.A(_3213_),
    .B(_3248_),
    .COUT(_3249_),
    .SUM(_3250_));
 sky130_fd_sc_hd__ha_1 _6905_ (.A(_3213_),
    .B(_3251_),
    .COUT(_3252_),
    .SUM(_3253_));
 sky130_fd_sc_hd__ha_4 _6906_ (.A(_3254_),
    .B(_3235_),
    .COUT(_3255_),
    .SUM(_3256_));
 sky130_fd_sc_hd__ha_1 _6907_ (.A(_3257_),
    .B(_3258_),
    .COUT(_3259_),
    .SUM(_3260_));
 sky130_fd_sc_hd__ha_1 _6908_ (.A(_3261_),
    .B(_3262_),
    .COUT(_3263_),
    .SUM(_3264_));
 sky130_fd_sc_hd__ha_1 _6909_ (.A(_3265_),
    .B(_3266_),
    .COUT(_3267_),
    .SUM(_3268_));
 sky130_fd_sc_hd__ha_1 _6910_ (.A(_3269_),
    .B(_3270_),
    .COUT(_3271_),
    .SUM(_3272_));
 sky130_fd_sc_hd__ha_1 _6911_ (.A(_3273_),
    .B(_3274_),
    .COUT(_3275_),
    .SUM(_3276_));
 sky130_fd_sc_hd__ha_1 _6912_ (.A(_3277_),
    .B(_3278_),
    .COUT(_3279_),
    .SUM(_3280_));
 sky130_fd_sc_hd__ha_1 _6913_ (.A(_3281_),
    .B(_3282_),
    .COUT(_3283_),
    .SUM(_3284_));
 sky130_fd_sc_hd__ha_1 _6914_ (.A(_3285_),
    .B(_3286_),
    .COUT(_3287_),
    .SUM(_3288_));
 sky130_fd_sc_hd__ha_1 _6915_ (.A(_2167_),
    .B(_2159_),
    .COUT(_3289_),
    .SUM(_3290_));
 sky130_fd_sc_hd__ha_1 _6916_ (.A(_3114_),
    .B(_3172_),
    .COUT(_2156_),
    .SUM(_3291_));
 sky130_fd_sc_hd__ha_1 _6917_ (.A(_3292_),
    .B(_3116_),
    .COUT(_2176_),
    .SUM(_3293_));
 sky130_fd_sc_hd__ha_2 _6918_ (.A(_3294_),
    .B(_3295_),
    .COUT(_3296_),
    .SUM(_3297_));
 sky130_fd_sc_hd__ha_1 _6919_ (.A(_3298_),
    .B(_3299_),
    .COUT(_3300_),
    .SUM(_3301_));
 sky130_fd_sc_hd__ha_1 _6920_ (.A(_3302_),
    .B(_3303_),
    .COUT(_3304_),
    .SUM(_3305_));
 sky130_fd_sc_hd__ha_1 _6921_ (.A(_3306_),
    .B(_3307_),
    .COUT(_3308_),
    .SUM(_3309_));
 sky130_fd_sc_hd__ha_2 _6922_ (.A(_3310_),
    .B(_3311_),
    .COUT(_3312_),
    .SUM(_3313_));
 sky130_fd_sc_hd__ha_1 _6923_ (.A(_3298_),
    .B(_3299_),
    .COUT(_3314_),
    .SUM(_3315_));
 sky130_fd_sc_hd__ha_2 _6924_ (.A(_3316_),
    .B(_3317_),
    .COUT(_3318_),
    .SUM(_3319_));
 sky130_fd_sc_hd__ha_1 _6925_ (.A(_3320_),
    .B(_3321_),
    .COUT(_3322_),
    .SUM(_3323_));
 sky130_fd_sc_hd__ha_1 _6926_ (.A(_3324_),
    .B(_3325_),
    .COUT(_3326_),
    .SUM(_3327_));
 sky130_fd_sc_hd__ha_2 _6927_ (.A(_3328_),
    .B(_3329_),
    .COUT(_3330_),
    .SUM(_3331_));
 sky130_fd_sc_hd__ha_1 _6928_ (.A(_3332_),
    .B(_3333_),
    .COUT(_3334_),
    .SUM(_3335_));
 sky130_fd_sc_hd__ha_1 _6929_ (.A(_3332_),
    .B(_3333_),
    .COUT(_3336_),
    .SUM(_3337_));
 sky130_fd_sc_hd__ha_1 _6930_ (.A(_3338_),
    .B(_3339_),
    .COUT(_3340_),
    .SUM(_3341_));
 sky130_fd_sc_hd__ha_1 _6931_ (.A(_3342_),
    .B(_3343_),
    .COUT(_3344_),
    .SUM(_3345_));
 sky130_fd_sc_hd__ha_1 _6932_ (.A(_3346_),
    .B(_3347_),
    .COUT(_3348_),
    .SUM(_3349_));
 sky130_fd_sc_hd__ha_1 _6933_ (.A(_3350_),
    .B(_3351_),
    .COUT(_3352_),
    .SUM(_3353_));
 sky130_fd_sc_hd__ha_1 _6934_ (.A(_3354_),
    .B(_3355_),
    .COUT(_3356_),
    .SUM(_3357_));
 sky130_fd_sc_hd__ha_1 _6935_ (.A(_2164_),
    .B(_2171_),
    .COUT(_3358_),
    .SUM(_3359_));
 sky130_fd_sc_hd__ha_1 _6936_ (.A(_3360_),
    .B(_3361_),
    .COUT(_3362_),
    .SUM(_3363_));
 sky130_fd_sc_hd__ha_1 _6937_ (.A(_3364_),
    .B(_3365_),
    .COUT(_3366_),
    .SUM(_3367_));
 sky130_fd_sc_hd__ha_1 _6938_ (.A(_3368_),
    .B(_3369_),
    .COUT(_3370_),
    .SUM(_3371_));
 sky130_fd_sc_hd__ha_2 _6939_ (.A(_3372_),
    .B(_3373_),
    .COUT(_3374_),
    .SUM(_3375_));
 sky130_fd_sc_hd__ha_1 _6940_ (.A(_3376_),
    .B(_3377_),
    .COUT(_3378_),
    .SUM(_3379_));
 sky130_fd_sc_hd__ha_1 _6941_ (.A(net7),
    .B(_3381_),
    .COUT(_3382_),
    .SUM(_3383_));
 sky130_fd_sc_hd__ha_1 _6942_ (.A(net7),
    .B(_3384_),
    .COUT(_3385_),
    .SUM(_3386_));
 sky130_fd_sc_hd__ha_1 _6943_ (.A(net7),
    .B(_3387_),
    .COUT(_3388_),
    .SUM(_3389_));
 sky130_fd_sc_hd__ha_1 _6944_ (.A(net7),
    .B(_3390_),
    .COUT(_3391_),
    .SUM(_3392_));
 sky130_fd_sc_hd__ha_1 _6945_ (.A(net7),
    .B(_3393_),
    .COUT(_3394_),
    .SUM(_3395_));
 sky130_fd_sc_hd__ha_1 _6946_ (.A(net7),
    .B(_3396_),
    .COUT(_3397_),
    .SUM(_3398_));
 sky130_fd_sc_hd__ha_1 _6947_ (.A(net7),
    .B(_3399_),
    .COUT(_3400_),
    .SUM(_3401_));
 sky130_fd_sc_hd__ha_1 _6948_ (.A(net20),
    .B(_3402_),
    .COUT(_3403_),
    .SUM(_3404_));
 sky130_fd_sc_hd__ha_1 _6949_ (.A(net8),
    .B(_3406_),
    .COUT(_3407_),
    .SUM(_3408_));
 sky130_fd_sc_hd__ha_1 _6950_ (.A(net20),
    .B(_3409_),
    .COUT(_3410_),
    .SUM(_3411_));
 sky130_fd_sc_hd__ha_1 _6951_ (.A(_3405_),
    .B(_3412_),
    .COUT(_3413_),
    .SUM(_3414_));
 sky130_fd_sc_hd__ha_1 _6952_ (.A(_3380_),
    .B(_3415_),
    .COUT(_3416_),
    .SUM(_3417_));
 sky130_fd_sc_hd__ha_1 _6953_ (.A(_3380_),
    .B(_3418_),
    .COUT(_3419_),
    .SUM(_3420_));
 sky130_fd_sc_hd__ha_4 _6954_ (.A(_3380_),
    .B(_3421_),
    .COUT(_3422_),
    .SUM(_3423_));
 sky130_fd_sc_hd__ha_2 _6955_ (.A(_3424_),
    .B(_3425_),
    .COUT(_3426_),
    .SUM(_3427_));
 sky130_fd_sc_hd__ha_1 _6956_ (.A(_3261_),
    .B(_3262_),
    .COUT(_3428_),
    .SUM(_3429_));
 sky130_fd_sc_hd__ha_1 _6957_ (.A(_3430_),
    .B(_3115_),
    .COUT(_3431_),
    .SUM(_3432_));
 sky130_fd_sc_hd__ha_1 _6958_ (.A(net178),
    .B(_3434_),
    .COUT(_3435_),
    .SUM(_3436_));
 sky130_fd_sc_hd__ha_2 _6959_ (.A(_3292_),
    .B(_3437_),
    .COUT(_3438_),
    .SUM(_3439_));
 sky130_fd_sc_hd__ha_4 _6960_ (.A(_3440_),
    .B(_3441_),
    .COUT(_3442_),
    .SUM(_3443_));
 sky130_fd_sc_hd__ha_1 _6961_ (.A(_3444_),
    .B(_3445_),
    .COUT(_3446_),
    .SUM(_3447_));
 sky130_fd_sc_hd__ha_1 _6962_ (.A(_3448_),
    .B(_3449_),
    .COUT(_3450_),
    .SUM(_3451_));
 sky130_fd_sc_hd__ha_1 _6963_ (.A(_3452_),
    .B(_3453_),
    .COUT(_3454_),
    .SUM(_3455_));
 sky130_fd_sc_hd__ha_1 _6964_ (.A(_2169_),
    .B(_2188_),
    .COUT(_3456_),
    .SUM(_3457_));
 sky130_fd_sc_hd__ha_1 _6965_ (.A(_3291_),
    .B(_3376_),
    .COUT(_2166_),
    .SUM(_3458_));
 sky130_fd_sc_hd__ha_1 _6966_ (.A(_3459_),
    .B(_3460_),
    .COUT(_3461_),
    .SUM(_3462_));
 sky130_fd_sc_hd__ha_1 _6967_ (.A(_2173_),
    .B(_2180_),
    .COUT(_3463_),
    .SUM(_3464_));
 sky130_fd_sc_hd__ha_1 _6968_ (.A(_3465_),
    .B(_3466_),
    .COUT(_3467_),
    .SUM(_3468_));
 sky130_fd_sc_hd__ha_2 _6969_ (.A(_3469_),
    .B(_3470_),
    .COUT(_3471_),
    .SUM(_3472_));
 sky130_fd_sc_hd__ha_1 _6970_ (.A(_3474_),
    .B(_3473_),
    .COUT(_3475_),
    .SUM(_3476_));
 sky130_fd_sc_hd__ha_1 _6971_ (.A(_3477_),
    .B(_3478_),
    .COUT(_3479_),
    .SUM(_3480_));
 sky130_fd_sc_hd__ha_1 _6972_ (.A(_3481_),
    .B(_3482_),
    .COUT(_3483_),
    .SUM(_3484_));
 sky130_fd_sc_hd__ha_2 _6973_ (.A(_3485_),
    .B(_3486_),
    .COUT(_3487_),
    .SUM(_3488_));
 sky130_fd_sc_hd__ha_1 _6974_ (.A(_3489_),
    .B(_3490_),
    .COUT(_3491_),
    .SUM(_3492_));
 sky130_fd_sc_hd__ha_1 _6975_ (.A(_3489_),
    .B(_3493_),
    .COUT(_3494_),
    .SUM(_3495_));
 sky130_fd_sc_hd__ha_1 _6976_ (.A(_3496_),
    .B(_3489_),
    .COUT(_3497_),
    .SUM(_3498_));
 sky130_fd_sc_hd__ha_1 _6977_ (.A(_3499_),
    .B(_3489_),
    .COUT(_3500_),
    .SUM(_3501_));
 sky130_fd_sc_hd__ha_1 _6978_ (.A(_3489_),
    .B(_3502_),
    .COUT(_3503_),
    .SUM(_3504_));
 sky130_fd_sc_hd__ha_1 _6979_ (.A(_3489_),
    .B(_3505_),
    .COUT(_3506_),
    .SUM(_3507_));
 sky130_fd_sc_hd__ha_1 _6980_ (.A(_3489_),
    .B(_3508_),
    .COUT(_3509_),
    .SUM(_3510_));
 sky130_fd_sc_hd__ha_1 _6981_ (.A(_3489_),
    .B(_3511_),
    .COUT(_3512_),
    .SUM(_3513_));
 sky130_fd_sc_hd__ha_1 _6982_ (.A(_3489_),
    .B(_3514_),
    .COUT(_3515_),
    .SUM(_3516_));
 sky130_fd_sc_hd__ha_1 _6983_ (.A(_3517_),
    .B(_3518_),
    .COUT(_3519_),
    .SUM(_3520_));
 sky130_fd_sc_hd__ha_1 _6984_ (.A(_3521_),
    .B(_3489_),
    .COUT(_3522_),
    .SUM(_3523_));
 sky130_fd_sc_hd__ha_1 _6985_ (.A(_2185_),
    .B(_2186_),
    .COUT(_3524_),
    .SUM(_3525_));
 sky130_fd_sc_hd__ha_4 _6986_ (.A(_3526_),
    .B(_2184_),
    .COUT(_3527_),
    .SUM(_3528_));
 sky130_fd_sc_hd__ha_1 _6987_ (.A(_3530_),
    .B(_3529_),
    .COUT(_3531_),
    .SUM(_3532_));
 sky130_fd_sc_hd__ha_1 _6988_ (.A(_3533_),
    .B(_3534_),
    .COUT(_3535_),
    .SUM(_3536_));
 sky130_fd_sc_hd__ha_1 _6989_ (.A(_3537_),
    .B(_3538_),
    .COUT(_3539_),
    .SUM(_3540_));
 sky130_fd_sc_hd__ha_1 _6990_ (.A(_3542_),
    .B(_3541_),
    .COUT(_3543_),
    .SUM(_3544_));
 sky130_fd_sc_hd__ha_1 _6991_ (.A(_3545_),
    .B(_3546_),
    .COUT(_3547_),
    .SUM(_3548_));
 sky130_fd_sc_hd__ha_1 _6992_ (.A(_3549_),
    .B(_3550_),
    .COUT(_3551_),
    .SUM(_3552_));
 sky130_fd_sc_hd__ha_2 _6993_ (.A(_3553_),
    .B(_3554_),
    .COUT(_3555_),
    .SUM(_3556_));
 sky130_fd_sc_hd__ha_1 _6994_ (.A(_3558_),
    .B(_3557_),
    .COUT(_3559_),
    .SUM(_3560_));
 sky130_fd_sc_hd__ha_1 _6995_ (.A(_3561_),
    .B(_3562_),
    .COUT(_3563_),
    .SUM(_3564_));
 sky130_fd_sc_hd__ha_2 _6996_ (.A(_3565_),
    .B(_3566_),
    .COUT(_3567_),
    .SUM(_3568_));
 sky130_fd_sc_hd__ha_2 _6997_ (.A(_3569_),
    .B(_3570_),
    .COUT(_3571_),
    .SUM(_3572_));
 sky130_fd_sc_hd__ha_1 _6998_ (.A(_3573_),
    .B(_3574_),
    .COUT(_3575_),
    .SUM(_3576_));
 sky130_fd_sc_hd__ha_1 _6999_ (.A(_3577_),
    .B(_3578_),
    .COUT(_3579_),
    .SUM(_3580_));
 sky130_fd_sc_hd__ha_2 _7000_ (.A(_3581_),
    .B(_3582_),
    .COUT(_3583_),
    .SUM(_3584_));
 sky130_fd_sc_hd__ha_2 _7001_ (.A(_3585_),
    .B(_3586_),
    .COUT(_3587_),
    .SUM(_3588_));
 sky130_fd_sc_hd__ha_1 _7002_ (.A(_3589_),
    .B(_3590_),
    .COUT(_3591_),
    .SUM(_3592_));
 sky130_fd_sc_hd__ha_1 _7003_ (.A(_3593_),
    .B(_3594_),
    .COUT(_3595_),
    .SUM(_3596_));
 sky130_fd_sc_hd__ha_4 _7004_ (.A(_3597_),
    .B(_3598_),
    .COUT(_3599_),
    .SUM(_3600_));
 sky130_fd_sc_hd__ha_1 _7005_ (.A(_3601_),
    .B(_3602_),
    .COUT(_3603_),
    .SUM(_3604_));
 sky130_fd_sc_hd__ha_4 _7006_ (.A(_3606_),
    .B(_3605_),
    .COUT(_3607_),
    .SUM(_3608_));
 sky130_fd_sc_hd__ha_4 _7007_ (.A(_3609_),
    .B(_3610_),
    .COUT(_3611_),
    .SUM(_3612_));
 sky130_fd_sc_hd__ha_1 _7008_ (.A(_3598_),
    .B(_3613_),
    .COUT(_3614_),
    .SUM(_3615_));
 sky130_fd_sc_hd__ha_1 _7009_ (.A(_3617_),
    .B(_3616_),
    .COUT(_3618_),
    .SUM(_3619_));
 sky130_fd_sc_hd__ha_1 _7010_ (.A(_3621_),
    .B(_3620_),
    .COUT(_3622_),
    .SUM(_3623_));
 sky130_fd_sc_hd__ha_1 _7011_ (.A(_3624_),
    .B(_3625_),
    .COUT(_3626_),
    .SUM(_3627_));
 sky130_fd_sc_hd__ha_1 _7012_ (.A(_3628_),
    .B(net154),
    .COUT(_3630_),
    .SUM(_3631_));
 sky130_fd_sc_hd__ha_1 _7013_ (.A(_3632_),
    .B(_3633_),
    .COUT(_3634_),
    .SUM(_3635_));
 sky130_fd_sc_hd__ha_1 _7014_ (.A(net134),
    .B(_3637_),
    .COUT(_3638_),
    .SUM(_3639_));
 sky130_fd_sc_hd__ha_2 _7015_ (.A(_3640_),
    .B(_3641_),
    .COUT(_3642_),
    .SUM(_3643_));
 sky130_fd_sc_hd__ha_1 _7016_ (.A(_3644_),
    .B(_3645_),
    .COUT(_3646_),
    .SUM(_3647_));
 sky130_fd_sc_hd__ha_2 _7017_ (.A(_3648_),
    .B(_3649_),
    .COUT(_3650_),
    .SUM(_3651_));
 sky130_fd_sc_hd__ha_1 _7018_ (.A(_3652_),
    .B(_3653_),
    .COUT(_3654_),
    .SUM(_3655_));
 sky130_fd_sc_hd__ha_2 _7019_ (.A(_3656_),
    .B(_3657_),
    .COUT(_3658_),
    .SUM(_3659_));
 sky130_fd_sc_hd__ha_1 _7020_ (.A(_3660_),
    .B(net224),
    .COUT(_3662_),
    .SUM(_3663_));
 sky130_fd_sc_hd__ha_2 _7021_ (.A(_3664_),
    .B(_3665_),
    .COUT(_3666_),
    .SUM(_3667_));
 sky130_fd_sc_hd__ha_1 _7022_ (.A(_3668_),
    .B(_3669_),
    .COUT(_3670_),
    .SUM(_3671_));
 sky130_fd_sc_hd__ha_4 _7023_ (.A(_3673_),
    .B(_3672_),
    .COUT(_3674_),
    .SUM(_3675_));
 sky130_fd_sc_hd__ha_4 _7024_ (.A(_2190_),
    .B(_2192_),
    .COUT(_3676_),
    .SUM(_3677_));
 sky130_fd_sc_hd__ha_1 _7025_ (.A(_3620_),
    .B(_3458_),
    .COUT(_2187_),
    .SUM(_3678_));
 sky130_fd_sc_hd__ha_4 _7026_ (.A(_3678_),
    .B(_3629_),
    .COUT(_2191_),
    .SUM(net78));
 sky130_fd_sc_hd__ha_4 _7027_ (.A(_3679_),
    .B(_3680_),
    .COUT(_3681_),
    .SUM(_3682_));
 sky130_fd_sc_hd__ha_2 _7028_ (.A(_3683_),
    .B(_3684_),
    .COUT(_3685_),
    .SUM(_3686_));
 sky130_fd_sc_hd__ha_4 _7029_ (.A(net67),
    .B(net68),
    .COUT(_3687_),
    .SUM(_3688_));
 sky130_fd_sc_hd__ha_4 _7030_ (.A(_3689_),
    .B(_3690_),
    .COUT(_3691_),
    .SUM(_3692_));
 sky130_fd_sc_hd__ha_1 _7031_ (.A(_3694_),
    .B(_3693_),
    .COUT(_3695_),
    .SUM(_3696_));
 sky130_fd_sc_hd__ha_1 _7032_ (.A(_3697_),
    .B(_3698_),
    .COUT(_3699_),
    .SUM(_3700_));
 sky130_fd_sc_hd__ha_1 _7033_ (.A(_3701_),
    .B(_3702_),
    .COUT(_3703_),
    .SUM(_3704_));
 sky130_fd_sc_hd__ha_4 _7034_ (.A(_3705_),
    .B(_3706_),
    .COUT(_3707_),
    .SUM(_3708_));
 sky130_fd_sc_hd__ha_1 _7035_ (.A(_3710_),
    .B(_3709_),
    .COUT(_3711_),
    .SUM(_3712_));
 sky130_fd_sc_hd__ha_1 _7036_ (.A(_3705_),
    .B(_3713_),
    .COUT(_3714_),
    .SUM(_3715_));
 sky130_fd_sc_hd__ha_1 _7037_ (.A(_3716_),
    .B(_3717_),
    .COUT(_3718_),
    .SUM(_3719_));
 sky130_fd_sc_hd__ha_4 _7038_ (.A(_3720_),
    .B(_3721_),
    .COUT(_3722_),
    .SUM(_3723_));
 sky130_fd_sc_hd__ha_1 _7039_ (.A(_3724_),
    .B(_3725_),
    .COUT(_3726_),
    .SUM(_3727_));
 sky130_fd_sc_hd__ha_1 _7040_ (.A(net118),
    .B(_3729_),
    .COUT(_3730_),
    .SUM(_3731_));
 sky130_fd_sc_hd__ha_1 _7041_ (.A(net138),
    .B(_3733_),
    .COUT(_3734_),
    .SUM(_3735_));
 sky130_fd_sc_hd__ha_1 _7042_ (.A(_3736_),
    .B(_3721_),
    .COUT(_3737_),
    .SUM(_3738_));
 sky130_fd_sc_hd__ha_1 _7043_ (.A(_3739_),
    .B(_3740_),
    .COUT(_3741_),
    .SUM(_3742_));
 sky130_fd_sc_hd__ha_1 _7044_ (.A(_3743_),
    .B(_3744_),
    .COUT(_3745_),
    .SUM(_3746_));
 sky130_fd_sc_hd__ha_4 _7045_ (.A(_3293_),
    .B(_3724_),
    .COUT(_2181_),
    .SUM(_3526_));
 sky130_fd_sc_hd__clkinv_2 clone1 (.A(_0629_),
    .Y(net1));
 sky130_fd_sc_hd__clkinv_2 clone3 (.A(_0158_),
    .Y(net3));
 sky130_fd_sc_hd__clkbuf_2 clone4 (.A(net5),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 split5 (.A(_2092_),
    .X(net5));
 sky130_fd_sc_hd__o21bai_4 clone6 (.A1(_0343_),
    .A2(_0342_),
    .B1_N(_0347_),
    .Y(net6));
 sky130_fd_sc_hd__clkbuf_4 clone7 (.A(_1185_),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 clone8 (.A(_1186_),
    .X(net8));
 sky130_fd_sc_hd__buf_6 clone9 (.A(net174),
    .X(net9));
 sky130_fd_sc_hd__buf_6 clone10 (.A(_1048_),
    .X(net10));
 sky130_fd_sc_hd__buf_6 clone11 (.A(_1049_),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 clone12 (.A(_0629_),
    .X(net12));
 sky130_fd_sc_hd__a311o_4 clone13 (.A1(_2660_),
    .A2(_0627_),
    .A3(_0626_),
    .B1(_0628_),
    .C1(_2653_),
    .X(net13));
 sky130_fd_sc_hd__buf_4 clone14 (.A(net174),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 clone15 (.A(_0159_),
    .X(net15));
 sky130_fd_sc_hd__clkinv_4 clone16 (.A(_0045_),
    .Y(net16));
 sky130_fd_sc_hd__clkbuf_2 clone17 (.A(_0873_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 clone18 (.A(_0158_),
    .X(net18));
 sky130_fd_sc_hd__buf_4 clone19 (.A(_1048_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 clone20 (.A(_1185_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 clone21 (.A(net211),
    .X(net21));
 sky130_fd_sc_hd__nand2b_2 clone22 (.A_N(_3382_),
    .B(_1315_),
    .Y(net22));
 sky130_fd_sc_hd__buf_4 clone23 (.A(_0295_),
    .X(net23));
 sky130_fd_sc_hd__buf_6 clone24 (.A(_0972_),
    .X(net24));
 sky130_fd_sc_hd__clkinv_4 clone25 (.A(_3213_),
    .Y(net25));
 sky130_fd_sc_hd__buf_4 clone26 (.A(_0972_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 clone27 (.A(_1319_),
    .X(net27));
 sky130_fd_sc_hd__buf_4 clone28 (.A(net62),
    .X(net28));
 sky130_fd_sc_hd__nor2_4 clone29 (.A(net205),
    .B(net202),
    .Y(net29));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(x_in[0]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(x_in[10]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(x_in[11]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(x_in[12]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(x_in[13]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(x_in[14]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(x_in[15]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(x_in[1]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(x_in[2]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(x_in[3]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(x_in[4]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(x_in[5]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(x_in[6]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(x_in[7]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(x_in[8]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(x_in[9]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(y_in[0]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(y_in[10]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(y_in[11]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(y_in[12]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(y_in[13]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(y_in[14]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(y_in[15]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(y_in[1]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(y_in[2]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(y_in[3]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(y_in[4]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(y_in[5]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(y_in[6]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(y_in[7]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(y_in[8]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(y_in[9]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input33 (.A(z_in[0]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(z_in[10]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(z_in[11]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(z_in[12]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(z_in[13]),
    .X(net66));
 sky130_fd_sc_hd__buf_8 input38 (.A(z_in[14]),
    .X(net67));
 sky130_fd_sc_hd__buf_6 input39 (.A(z_in[15]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(z_in[1]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(z_in[2]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(z_in[3]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(z_in[4]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(z_in[5]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(z_in[6]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(z_in[7]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(z_in[8]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(z_in[9]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net78),
    .X(x_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net79),
    .X(x_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net80),
    .X(x_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net81),
    .X(x_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net82),
    .X(x_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net83),
    .X(x_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net84),
    .X(x_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net85),
    .X(x_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net86),
    .X(x_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net87),
    .X(x_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net88),
    .X(x_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net89),
    .X(x_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net90),
    .X(x_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net91),
    .X(x_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net92),
    .X(x_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net93),
    .X(x_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net94),
    .X(y_out[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net95),
    .X(y_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net96),
    .X(y_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net97),
    .X(y_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net98),
    .X(y_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net99),
    .X(y_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net100),
    .X(y_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net101),
    .X(y_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net102),
    .X(y_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net103),
    .X(y_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net104),
    .X(y_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net105),
    .X(y_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net106),
    .X(y_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net107),
    .X(y_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net108),
    .X(y_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net109),
    .X(y_out[9]));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(_1545_),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer2 (.A(net200),
    .X(net111));
 sky130_fd_sc_hd__buf_6 rebuffer3 (.A(net111),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_3264_),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_1223_),
    .X(net114));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(_3476_),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net115),
    .X(net116));
 sky130_fd_sc_hd__buf_4 rebuffer8 (.A(_1351_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net158),
    .X(net118));
 sky130_fd_sc_hd__buf_2 rebuffer10 (.A(_1965_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 rebuffer11 (.A(_2000_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net205),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(_1413_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(_1328_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net123),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(net123),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer17 (.A(net125),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(_1401_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(_1221_),
    .X(net128));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(_2193_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(_1289_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(_1510_),
    .X(net131));
 sky130_fd_sc_hd__buf_6 rebuffer78 (.A(_1564_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(_3532_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(_3636_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net148),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(_1326_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(_3732_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(_3732_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(_1121_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(_1291_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(_1427_),
    .X(net141));
 sky130_fd_sc_hd__buf_6 rebuffer33 (.A(_1994_),
    .X(net142));
 sky130_fd_sc_hd__buf_4 rebuffer34 (.A(net207),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 rebuffer35 (.A(_3544_),
    .X(net144));
 sky130_fd_sc_hd__buf_6 rebuffer36 (.A(_1501_),
    .X(net145));
 sky130_fd_sc_hd__buf_4 rebuffer37 (.A(_1532_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net211),
    .X(net147));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer39 (.A(_1329_),
    .X(net148));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer40 (.A(net212),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(_1512_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(_1514_),
    .X(net151));
 sky130_fd_sc_hd__buf_4 rebuffer43 (.A(_2006_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(_3629_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net153),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(_1495_),
    .X(net155));
 sky130_fd_sc_hd__buf_2 rebuffer47 (.A(_1340_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 rebuffer48 (.A(_3728_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net157),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net214),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(_1293_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_1 rebuffer61 (.A(_1369_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_16 clone62 (.A(_0008_),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_16 clone63 (.A(_0010_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_16 clone67 (.A(_0009_),
    .X(net176));
 sky130_fd_sc_hd__buf_6 rebuffer68 (.A(_1327_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(_3433_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(net178),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer79 (.A(_1472_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(_1469_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 rebuffer81 (.A(_1535_),
    .X(net190));
 sky130_fd_sc_hd__buf_6 rebuffer82 (.A(_1535_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(_3606_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net192),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(_1205_),
    .X(net194));
 sky130_fd_sc_hd__buf_2 rebuffer112 (.A(_1929_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer113 (.A(_1499_),
    .X(net222));
 sky130_fd_sc_hd__buf_6 rebuffer114 (.A(_1529_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer115 (.A(_3661_),
    .X(net224));
 sky130_fd_sc_hd__buf_2 rebuffer119 (.A(_1925_),
    .X(net228));
 sky130_fd_sc_hd__buf_2 rebuffer120 (.A(_1936_),
    .X(net229));
 sky130_fd_sc_hd__buf_6 rebuffer124 (.A(_1927_),
    .X(net233));
 sky130_fd_sc_hd__buf_2 rebuffer126 (.A(_1940_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 rebuffer127 (.A(net235),
    .X(net236));
 sky130_fd_sc_hd__buf_1 rebuffer128 (.A(_1516_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 rebuffer129 (.A(_3672_),
    .X(net238));
 sky130_fd_sc_hd__buf_6 rebuffer130 (.A(_2194_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 rebuffer131 (.A(_2183_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 rebuffer132 (.A(_2021_),
    .X(net241));
 sky130_fd_sc_hd__buf_1 rebuffer133 (.A(net241),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(_3560_),
    .X(net173));
 sky130_fd_sc_hd__buf_4 rebuffer63 (.A(_0348_),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer64 (.A(_1376_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(_1504_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net180),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer76 (.A(_1491_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(_1969_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer86 (.A(net197),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer87 (.A(net205),
    .X(net199));
 sky130_fd_sc_hd__buf_1 rebuffer88 (.A(_1545_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer89 (.A(_3706_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer90 (.A(_1469_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(net202),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer92 (.A(net202),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer93 (.A(_1470_),
    .X(net205));
 sky130_fd_sc_hd__buf_1 rebuffer94 (.A(_1528_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 rebuffer95 (.A(_1531_),
    .X(net207));
 sky130_fd_sc_hd__buf_2 rebuffer96 (.A(_1917_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 rebuffer97 (.A(_3696_),
    .X(net209));
 sky130_fd_sc_hd__buf_2 rebuffer98 (.A(_1935_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer99 (.A(_1318_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer100 (.A(net211),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer101 (.A(_3623_),
    .X(net213));
 sky130_fd_sc_hd__buf_2 rebuffer102 (.A(_3728_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 rebuffer103 (.A(_2018_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer152 (.A(_1273_),
    .X(net264));
 sky130_fd_sc_hd__buf_1 rebuffer160 (.A(_1520_),
    .X(net272));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
endmodule
